// Copyright 2023 Flavien Solt, ETH Zurich.
// Licensed under the General Public License, Version 3.0, see LICENSE for details.
// SPDX-License-Identifier: GPL-3.0-only

module top(in_data, out_data);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  reg _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  reg _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  reg _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  reg _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  reg _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire [16:0] _1886_;
  wire [16:0] _1887_;
  wire [13:0] _1888_;
  wire [12:0] _1889_;
  wire [12:0] _1890_;
  wire [12:0] _1891_;
  wire [55:0] _1892_;
  wire [55:0] _1893_;
  wire [55:0] _1894_;
  wire [35:0] _1895_;
  wire [35:0] _1896_;
  wire [53:0] _1897_;
  wire [53:0] _1898_;
  wire [53:0] _1899_;
  wire [86:0] _1900_;
  wire [86:0] _1901_;
  wire [38:0] _1902_;
  wire [38:0] _1903_;
  wire [38:0] _1904_;
  wire [4:0] _1905_;
  wire [4:0] _1906_;
  wire [55:0] _1907_;
  wire [39:0] _1908_;
  wire [39:0] _1909_;
  wire [9:0] _1910_;
  wire [14:0] _1911_;
  wire [39:0] _1912_;
  wire [39:0] _1913_;
  wire [46:0] _1914_;
  wire [46:0] _1915_;
  wire [8:0] _1916_;
  wire [13:0] _1917_;
  wire [31:0] _1918_;
  wire [31:0] _1919_;
  wire [31:0] _1920_;
  wire _1921_;
  wire [2:0] _1922_;
  wire [7:0] _1923_;
  wire [7:0] _1924_;
  wire [30:0] _1925_;
  wire [30:0] _1926_;
  wire [24:0] _1927_;
  wire [24:0] _1928_;
  wire [27:0] _1929_;
  wire [27:0] _1930_;
  wire [3:0] _1931_;
  wire [12:0] _1932_;
  wire [29:0] _1933_;
  wire [5:0] _1934_;
  wire [79:0] _1935_;
  wire [79:0] _1936_;
  wire [1:0] _1937_;
  wire [8:0] _1938_;
  wire [12:0] _1939_;
  wire [37:0] _1940_;
  wire [37:0] _1941_;
  wire [111:0] _1942_;
  wire [111:0] _1943_;
  wire [35:0] _1944_;
  wire [7:0] _1945_;
  wire [13:0] _1946_;
  wire [13:0] _1947_;
  wire [9:0] _1948_;
  wire [9:0] _1949_;
  wire [215:0] _1950_;
  wire [215:0] _1951_;
  wire [215:0] _1952_;
  wire [28:0] _1953_;
  wire [28:0] _1954_;
  wire [30:0] _1955_;
  wire [30:0] _1956_;
  wire [13:0] _1957_;
  wire [13:0] _1958_;
  wire [9:0] _1959_;
  wire [34:0] _1960_;
  wire [34:0] _1961_;
  wire [34:0] _1962_;
  wire [76:0] _1963_;
  wire [76:0] _1964_;
  wire [77:0] _1965_;
  wire [77:0] _1966_;
  wire [77:0] _1967_;
  wire [51:0] _1968_;
  wire [51:0] _1969_;
  wire [51:0] _1970_;
  wire [25:0] _1971_;
  wire [25:0] _1972_;
  wire [25:0] _1973_;
  wire [1:0] _1974_;
  wire [74:0] _1975_;
  wire [74:0] _1976_;
  wire [74:0] _1977_;
  wire [58:0] _1978_;
  wire [58:0] _1979_;
  wire [23:0] _1980_;
  wire [23:0] _1981_;
  wire [23:0] _1982_;
  wire [46:0] _1983_;
  wire [46:0] _1984_;
  wire [11:0] _1985_;
  wire [11:0] _1986_;
  wire [54:0] _1987_;
  wire [54:0] _1988_;
  wire [54:0] _1989_;
  wire [55:0] _1990_;
  wire [55:0] _1991_;
  wire [55:0] _1992_;
  wire [9:0] _1993_;
  wire [9:0] _1994_;
  wire [17:0] _1995_;
  wire [17:0] _1996_;
  wire [2:0] _1997_;
  wire [40:0] _1998_;
  wire [139:0] _1999_;
  wire [139:0] _2000_;
  wire [139:0] _2001_;
  wire [31:0] _2002_;
  wire [10:0] _2003_;
  wire [10:0] _2004_;
  wire [10:0] _2005_;
  wire [8:0] _2006_;
  wire [8:0] _2007_;
  wire [14:0] _2008_;
  wire [3:0] _2009_;
  wire [3:0] _2010_;
  wire [43:0] _2011_;
  wire [43:0] _2012_;
  wire [17:0] _2013_;
  wire [17:0] _2014_;
  wire [21:0] _2015_;
  wire [21:0] _2016_;
  wire [65:0] _2017_;
  wire [65:0] _2018_;
  wire [65:0] _2019_;
  wire [27:0] _2020_;
  wire [21:0] _2021_;
  wire [21:0] _2022_;
  wire [13:0] _2023_;
  wire [13:0] _2024_;
  wire [43:0] _2025_;
  wire [43:0] _2026_;
  wire [10:0] _2027_;
  wire [10:0] _2028_;
  wire [43:0] _2029_;
  wire [66:0] _2030_;
  wire [66:0] _2031_;
  wire [66:0] _2032_;
  wire [23:0] _2033_;
  wire [23:0] _2034_;
  wire [23:0] _2035_;
  wire [16:0] _2036_;
  wire [80:0] _2037_;
  wire [80:0] _2038_;
  wire [13:0] _2039_;
  wire [35:0] _2040_;
  wire [35:0] _2041_;
  wire [12:0] _2042_;
  wire [12:0] _2043_;
  wire [8:0] _2044_;
  wire [8:0] _2045_;
  wire [21:0] _2046_;
  wire [83:0] _2047_;
  wire [83:0] _2048_;
  wire [83:0] _2049_;
  wire [9:0] _2050_;
  wire [9:0] _2051_;
  wire [40:0] _2052_;
  wire [40:0] _2053_;
  wire [40:0] _2054_;
  wire [3:0] _2055_;
  wire [3:0] _2056_;
  wire [2:0] _2057_;
  wire [95:0] _2058_;
  wire [95:0] _2059_;
  wire [95:0] _2060_;
  wire [10:0] _2061_;
  wire [43:0] _2062_;
  wire [43:0] _2063_;
  wire [43:0] _2064_;
  wire [57:0] _2065_;
  wire [9:0] _2066_;
  wire [5:0] _2067_;
  wire [32:0] _2068_;
  wire [32:0] _2069_;
  wire [32:0] _2070_;
  wire [44:0] _2071_;
  wire [44:0] _2072_;
  wire [6:0] _2073_;
  wire [6:0] _2074_;
  wire [14:0] _2075_;
  wire [28:0] _2076_;
  wire [20:0] _2077_;
  wire [21:0] _2078_;
  wire [21:0] _2079_;
  wire [31:0] _2080_;
  wire [31:0] _2081_;
  wire [31:0] _2082_;
  wire [28:0] _2083_;
  wire [9:0] _2084_;
  wire [9:0] _2085_;
  wire [31:0] _2086_;
  wire [31:0] _2087_;
  wire [22:0] _2088_;
  wire [5:0] _2089_;
  wire [14:0] _2090_;
  wire [14:0] _2091_;
  wire [14:0] _2092_;
  wire [130:0] _2093_;
  wire [130:0] _2094_;
  wire [130:0] _2095_;
  wire [39:0] _2096_;
  wire [39:0] _2097_;
  wire [39:0] _2098_;
  wire [9:0] _2099_;
  wire [165:0] _2100_;
  wire [165:0] _2101_;
  wire [165:0] _2102_;
  wire [6:0] _2103_;
  wire [6:0] _2104_;
  wire [43:0] _2105_;
  wire [30:0] _2106_;
  wire [30:0] _2107_;
  wire [84:0] _2108_;
  wire [8:0] _2109_;
  wire [51:0] _2110_;
  wire [51:0] _2111_;
  wire [97:0] _2112_;
  wire [25:0] _2113_;
  wire [25:0] _2114_;
  wire [14:0] _2115_;
  wire [8:0] _2116_;
  wire [8:0] _2117_;
  wire [99:0] _2118_;
  wire [99:0] _2119_;
  wire [99:0] _2120_;
  wire [97:0] _2121_;
  wire [22:0] _2122_;
  wire [22:0] _2123_;
  wire [14:0] _2124_;
  wire [48:0] _2125_;
  wire [48:0] _2126_;
  wire [6:0] _2127_;
  wire [16:0] _2128_;
  wire [16:0] _2129_;
  wire [6:0] _2130_;
  wire [1:0] _2131_;
  wire [1:0] _2132_;
  wire [6:0] _2133_;
  wire [6:0] _2134_;
  wire [7:0] _2135_;
  wire [8:0] _2136_;
  wire [2:0] _2137_;
  wire [72:0] _2138_;
  wire [72:0] _2139_;
  wire [22:0] _2140_;
  wire [22:0] _2141_;
  wire [84:0] _2142_;
  wire [84:0] _2143_;
  wire [63:0] _2144_;
  wire [23:0] _2145_;
  wire [23:0] _2146_;
  wire [5:0] _2147_;
  wire [60:0] _2148_;
  wire [60:0] _2149_;
  wire [60:0] _2150_;
  wire [34:0] _2151_;
  wire [3:0] _2152_;
  wire [39:0] _2153_;
  wire [39:0] _2154_;
  wire [11:0] _2155_;
  wire [102:0] _2156_;
  wire [38:0] _2157_;
  wire [50:0] _2158_;
  wire [50:0] _2159_;
  wire [50:0] _2160_;
  wire [28:0] _2161_;
  wire [42:0] _2162_;
  wire [42:0] _2163_;
  wire [29:0] _2164_;
  wire [46:0] _2165_;
  wire [46:0] _2166_;
  wire [6:0] _2167_;
  wire [169:0] _2168_;
  wire [169:0] _2169_;
  wire [169:0] _2170_;
  wire [2:0] _2171_;
  wire [23:0] _2172_;
  wire [23:0] _2173_;
  wire [9:0] _2174_;
  wire [12:0] _2175_;
  wire [7:0] _2176_;
  wire [33:0] _2177_;
  wire [81:0] _2178_;
  wire [6:0] _2179_;
  wire [6:0] _2180_;
  wire [11:0] _2181_;
  wire [102:0] _2182_;
  wire [102:0] _2183_;
  wire [13:0] _2184_;
  wire [64:0] _2185_;
  wire [28:0] _2186_;
  wire [24:0] _2187_;
  wire [24:0] _2188_;
  wire [78:0] _2189_;
  wire [78:0] _2190_;
  wire [9:0] _2191_;
  wire [37:0] _2192_;
  wire [7:0] _2193_;
  wire [10:0] _2194_;
  wire [10:0] _2195_;
  wire [154:0] _2196_;
  wire [154:0] _2197_;
  wire [47:0] _2198_;
  wire [47:0] _2199_;
  wire [47:0] _2200_;
  wire [12:0] _2201_;
  wire [4:0] _2202_;
  wire [17:0] _2203_;
  wire [2:0] _2204_;
  wire [19:0] _2205_;
  wire [11:0] _2206_;
  wire [4:0] _2207_;
  wire [3:0] _2208_;
  wire [32:0] _2209_;
  wire [13:0] _2210_;
  wire [13:0] _2211_;
  wire [6:0] _2212_;
  wire [23:0] _2213_;
  wire [23:0] _2214_;
  wire [7:0] _2215_;
  wire [100:0] _2216_;
  wire [43:0] _2217_;
  wire [43:0] _2218_;
  wire [43:0] _2219_;
  wire [82:0] _2220_;
  wire [82:0] _2221_;
  wire [1:0] _2222_;
  wire [55:0] _2223_;
  wire [17:0] _2224_;
  wire [64:0] _2225_;
  wire [67:0] _2226_;
  wire [38:0] _2227_;
  wire [67:0] _2228_;
  wire [67:0] _2229_;
  wire [12:0] _2230_;
  wire [197:0] _2231_;
  wire [7:0] _2232_;
  wire [52:0] _2233_;
  wire [32:0] _2234_;
  wire [66:0] _2235_;
  wire [66:0] _2236_;
  wire [40:0] _2237_;
  wire [122:0] _2238_;
  wire _2239_;
  wire [72:0] _2240_;
  wire [39:0] _2241_;
  wire [21:0] _2242_;
  wire [12:0] _2243_;
  wire [82:0] _2244_;
  wire [82:0] _2245_;
  wire [1:0] _2246_;
  wire _2247_;
  wire [35:0] _2248_;
  wire [40:0] _2249_;
  wire [70:0] _2250_;
  wire [16:0] _2251_;
  wire _2252_;
  wire [6:0] _2253_;
  wire [54:0] _2254_;
  wire [34:0] _2255_;
  wire [65:0] _2256_;
  wire [36:0] _2257_;
  wire [59:0] _2258_;
  wire [53:0] _2259_;
  wire [42:0] _2260_;
  wire [109:0] _2261_;
  wire [109:0] _2262_;
  wire [59:0] _2263_;
  wire [90:0] _2264_;
  wire [61:0] _2265_;
  wire [104:0] _2266_;
  wire [10:0] _2267_;
  wire [98:0] _2268_;
  wire [12:0] _2269_;
  wire [76:0] _2270_;
  wire [48:0] _2271_;
  wire [23:0] _2272_;
  wire [69:0] _2273_;
  wire [33:0] _2274_;
  reg [13:0] _2275_;
  wire [64:0] _2276_;
  wire _2277_;
  wire [56:0] _2278_;
  wire [55:0] _2279_;
  wire [64:0] _2280_;
  wire [82:0] _2281_;
  wire [119:0] _2282_;
  wire [120:0] _2283_;
  wire [40:0] _2284_;
  wire [81:0] _2285_;
  wire [14:0] _2286_;
  wire [29:0] _2287_;
  wire [4:0] _2288_;
  wire [121:0] _2289_;
  wire [52:0] _2290_;
  wire [23:0] _2291_;
  wire [1:0] _2292_;
  wire [14:0] _2293_;
  wire [13:0] _2294_;
  wire [31:0] _2295_;
  wire [10:0] _2296_;
  wire [24:0] _2297_;
  wire [29:0] _2298_;
  wire [26:0] _2299_;
  wire [24:0] _2300_;
  wire [24:0] _2301_;
  wire [55:0] _2302_;
  wire [60:0] _2303_;
  reg [2:0] _2304_;
  wire [26:0] _2305_;
  wire [43:0] _2306_;
  wire [29:0] _2307_;
  wire [104:0] _2308_;
  wire [12:0] _2309_;
  wire [61:0] _2310_;
  wire [55:0] _2311_;
  wire [1:0] _2312_;
  wire [30:0] _2313_;
  wire [29:0] _2314_;
  wire [133:0] _2315_;
  wire [6:0] _2316_;
  wire [46:0] _2317_;
  wire [14:0] _2318_;
  wire [167:0] _2319_;
  wire [14:0] _2320_;
  wire [52:0] _2321_;
  wire [68:0] _2322_;
  wire [33:0] _2323_;
  input [2271:0] in_data;
  wire [2271:0] in_data;
  output [2047:0] out_data;
  wire [2047:0] out_data;
  assign _0015_ = _0019_ & ~(_0018_);
  assign _0029_ = _0031_ & ~(_0030_);
  assign _0042_ = _0044_ & ~(_0043_);
  assign _0051_ = _0053_ & ~(_0052_);
  assign _0060_ = _0062_ & ~(_0061_);
  assign _0067_ = _0069_ & ~(_0068_);
  assign out_data[1664] = _0075_ & ~(_0074_);
  assign out_data[1568] = _0077_ & ~(_0076_);
  assign out_data[1536] = _0079_ & ~(_0078_);
  assign out_data[832] = _0083_ & ~(_0081_);
  assign _0080_ = _0084_ & ~(_0082_);
  assign out_data[704] = _0060_ & ~(_0085_);
  assign out_data[320] = _0087_ & ~(_0086_);
  assign out_data[192] = _0089_ & ~(_0088_);
  assign out_data[128] = _0091_ & ~(_0090_);
  assign _0092_ = _0094_ & ~(_0093_);
  assign _0095_ = _0097_ & ~(_0096_);
  assign _0098_ = _0100_ & ~(_0099_);
  assign _0102_ = _0018_ & ~(_0103_);
  assign _0068_ = _0104_ & ~(_0101_);
  assign _0105_ = _0107_ & ~(_0106_);
  assign _0108_ = _0096_ & ~(_0109_);
  assign _0110_ = _0111_ & ~(_0065_);
  assign _0112_ = _0114_ & ~(_0113_);
  assign _0115_ = _0116_ & ~(_0042_);
  assign _0117_ = _0059_ & ~(_0118_);
  assign _0119_ = _0121_ & ~(_0120_);
  assign _0122_ = _0124_ & ~(_0123_);
  assign _0125_ = _0127_ & ~(_0126_);
  assign _0129_ = _0131_ & ~(_0130_);
  assign _0133_ = _0134_ & ~(_0016_);
  assign _0135_ = _0136_ & ~(_0025_);
  assign _0128_ = _0134_ & ~(_0132_);
  assign _0137_ = _0139_ & ~(_0138_);
  assign _0140_ = _0142_ & ~(_0141_);
  assign _0143_ = _0144_ & ~(_0096_);
  assign _0145_ = _0147_ & ~(_0146_);
  assign _0148_ = _0151_ & ~(_0149_);
  assign _0153_ = _0122_ & ~(_0152_);
  assign _0150_ = _0125_ & ~(_0152_);
  assign _0052_ = _0155_ & ~(_0154_);
  assign _0041_ = _0157_ & ~(_0156_);
  assign _0158_ = _0160_ & ~(_0159_);
  assign _0161_ = _0025_ & ~(_0162_);
  assign _0062_ = _0140_ & ~(_0163_);
  assign _0164_ = _0025_ & ~(_0165_);
  assign _0166_ = _0167_ & ~(_0138_);
  assign _0168_ = _0169_ & ~(_0135_);
  assign _0170_ = _0172_ & ~(_0171_);
  assign _0173_ = _0175_ & ~(_0174_);
  assign _0176_ = _0178_ & ~(_0177_);
  assign _0179_ = _0181_ & ~(_0180_);
  assign _0182_ = _0166_ & ~(_0132_);
  assign _0183_ = _0132_ & ~(_0109_);
  assign _0184_ = _0186_ & ~(_0185_);
  assign _0187_ = _0134_ & ~(_0188_);
  assign _0190_ = _0049_ & ~(_0191_);
  assign _0192_ = _0194_ & ~(_0193_);
  assign _0195_ = _0197_ & ~(_0196_);
  assign _0053_ = _0152_ & ~(_0198_);
  assign _0199_ = _0200_ & ~(_0084_);
  assign _0201_ = _0195_ & ~(_0200_);
  assign _0202_ = _0204_ & ~(_0203_);
  assign _0189_ = _0101_ & ~(_0025_);
  assign _0205_ = _0206_ & ~(_0149_);
  assign _0207_ = _0032_ & ~(_0208_);
  assign _0209_ = _0210_ & ~(_0096_);
  assign out_data[896] = _0212_ & ~(_0211_);
  assign _0213_ = _0215_ & ~(_0214_);
  assign _0216_ = _0217_ & ~(_0068_);
  assign _0218_ = _0219_ & ~(_0194_);
  assign _0220_ = _0221_ & ~(_0046_);
  assign _0222_ = _0224_ & ~(_0223_);
  assign _0225_ = _0112_ & ~(_0226_);
  assign _0227_ = _0068_ & ~(_0228_);
  assign _0229_ = _0231_ & ~(_0230_);
  assign _0234_ = _0236_ & ~(_0235_);
  assign _0232_ = _0237_ & ~(_0233_);
  assign _0239_ = _0240_ & ~(_0015_);
  assign _0005_ = _0243_ & ~(_0242_);
  assign _0047_ = _0182_ & ~(_0244_);
  assign _0245_ = _0057_ & ~(_0246_);
  assign _0247_ = _0249_ & ~(_0248_);
  assign _0010_ = _0252_ & ~(_0251_);
  assign _0253_ = _0254_ & ~(_0096_);
  assign _0238_ = _0250_ & ~(_0241_);
  assign _0255_ = _0256_ & ~(_0013_);
  assign _0257_ = _0258_ & ~(_0043_);
  assign _0261_ = _0262_ & ~(_0014_);
  assign _0263_ = _0210_ & ~(_0264_);
  assign _0265_ = _0068_ & ~(_0084_);
  assign _0266_ = _0058_ & ~(_0267_);
  assign _0268_ = _0270_ & ~(_0269_);
  assign _0271_ = _0019_ & ~(_0272_);
  assign _0273_ = _0275_ & ~(_0274_);
  assign _0276_ = _0278_ & ~(_0277_);
  assign _0279_ = _0281_ & ~(_0280_);
  assign _0282_ = _0283_ & ~(_0194_);
  assign _0284_ = _0286_ & ~(_0285_);
  assign _0288_ = _0289_ & ~(_0140_);
  assign _0292_ = _0190_ & ~(_0293_);
  assign _0295_ = _0144_ & ~(_0296_);
  assign _0290_ = _0294_ & ~(_0291_);
  assign _0297_ = _0299_ & ~(_0298_);
  assign _0300_ = _0297_ & ~(_0301_);
  assign _0302_ = _0303_ & ~(_0193_);
  assign _0305_ = _0307_ & ~(_0306_);
  assign _0304_ = _0194_ & ~(_0097_);
  assign _0308_ = _0309_ & ~(_0190_);
  assign _0310_ = _0311_ & ~(_0133_);
  assign _0312_ = _0314_ & ~(_0313_);
  assign _0315_ = _0317_ & ~(_0316_);
  assign _0318_ = _0320_ & ~(_0319_);
  assign _0321_ = _0322_ & ~(_0281_);
  assign _0326_ = _0327_ & ~(out_data[416]);
  assign _0030_ = _0329_ & ~(_0328_);
  assign _0330_ = _0332_ & ~(_0331_);
  assign _0333_ = _0335_ & ~(_0334_);
  assign _0336_ = _0338_ & ~(_0337_);
  assign _0339_ = _0340_ & ~(_0121_);
  assign _0341_ = _0342_ & ~(_0214_);
  assign _0343_ = _0154_ & ~(_0344_);
  assign _0026_ = _0332_ & ~(_0345_);
  assign _0347_ = _0348_ & ~(_0325_);
  assign _0349_ = _0351_ & ~(_0350_);
  assign _0352_ = _0354_ & ~(_0353_);
  assign _0355_ = _0356_ & ~(_0016_);
  assign _0358_ = _0359_ & ~(_0119_);
  assign _0360_ = _0362_ & ~(_0361_);
  assign _0363_ = _0221_ & ~(_0364_);
  assign _0366_ = _0257_ & ~(_0333_);
  assign _0367_ = _0368_ & ~(_0018_);
  assign _0370_ = _0371_ & ~(_0036_);
  assign _0372_ = _0253_ & ~(_0373_);
  assign _0374_ = _0376_ & ~(_0375_);
  assign _0377_ = _0379_ & ~(_0378_);
  assign _0381_ = _0383_ & ~(_0382_);
  assign _0384_ = _0386_ & ~(_0385_);
  assign _0387_ = _0389_ & ~(_0388_);
  assign _0390_ = _0391_ & ~(_0061_);
  assign _0392_ = _0311_ & ~(_0168_);
  assign _0393_ = _0096_ & ~(_0394_);
  assign _0395_ = _0397_ & ~(_0396_);
  assign _0398_ = _0399_ & ~(_0019_);
  assign _0400_ = _0402_ & ~(_0401_);
  assign _0109_ = _0404_ & ~(_0227_);
  assign _0405_ = _0407_ & ~(_0406_);
  assign _0408_ = _0410_ & ~(_0409_);
  assign _0413_ = _0414_ & ~(_0229_);
  assign _0415_ = _0416_ & ~(_0395_);
  assign _0277_ = _0241_ & ~(in_data[492]);
  assign _0421_ = _0422_ & ~(_0286_);
  assign _0423_ = _0357_ & ~(_0424_);
  assign _0426_ = _0428_ & ~(_0427_);
  assign _0429_ = _0431_ & ~(_0430_);
  assign _0435_ = _0437_ & ~(_0436_);
  assign _0439_ = _0441_ & ~(_0440_);
  assign _0442_ = _0208_ & ~(_0443_);
  assign _0445_ = _0446_ & ~(_0355_);
  assign _0025_ = _0241_ & ~(_0241_);
  assign _0449_ = _0451_ & ~(_0450_);
  assign out_data[1888] = _0458_ & ~(_0457_);
  assign _0217_ = _0464_ & ~(_0463_);
  assign _0465_ = _0467_ & ~(_0466_);
  assign _0470_ = _0239_ & ~(_0471_);
  assign _0472_ = _0474_ & ~(_0473_);
  assign _0476_ = _0477_ & ~(_0451_);
  assign _0480_ = _0482_ & ~(_0481_);
  assign _0483_ = _0485_ & ~(_0484_);
  assign _0493_ = _0495_ & ~(_0494_);
  assign _0496_ = _0497_ & ~(_0018_);
  assign _0096_ = _0189_ & ~(_0499_);
  assign _0512_ = _0514_ & ~(_0513_);
  assign _0517_ = _0058_ & ~(_0518_);
  assign _0521_ = _0210_ & _0522_;
  assign _0526_ = _0528_ & _0527_;
  assign out_data[1024] = _0016_ & _0532_;
  assign _0533_ = _0535_ & _0534_;
  assign _0529_ = _0206_ & _0277_;
  assign _0542_ = _0544_ & _0543_;
  assign _0554_ = _0227_ & _0553_;
  assign _0563_ = _0565_ & _0564_;
  assign _0568_ = _0569_ & _0287_;
  assign _0566_ = _0096_ & _0134_;
  assign _0570_ = _0003_ & _0571_;
  assign _0572_ = _0316_ & _0573_;
  assign _0134_ = in_data[1039] & _0033_;
  assign out_data[1440] = _0578_ & _0515_;
  assign out_data[1056] = _0579_ & _0347_;
  assign out_data[672] = _0580_ & _0003_;
  assign out_data[640] = _0582_ & _0581_;
  assign out_data[384] = _0584_ & _0583_;
  assign out_data[96] = _0586_ & _0585_;
  assign _0274_ = _0529_ & _0311_;
  assign _0587_ = _0589_ & _0588_;
  assign _0590_ = _0097_ & _0591_;
  assign _0335_ = _0098_ & _0592_;
  assign _0593_ = _0250_ & _0438_;
  assign _0309_ = _0095_ & _0306_;
  assign _0038_ = _0189_ & _0082_;
  assign _0594_ = _0589_ & _0595_;
  assign _0243_ = _0057_ & _0217_;
  assign _0485_ = _0316_ & _0152_;
  assign _0259_ = _0597_ & _0596_;
  assign _0598_ = _0227_ & _0599_;
  assign _0324_ = _0071_ & _0134_;
  assign _0600_ = _0601_ & _0084_;
  assign _0419_ = _0603_ & _0602_;
  assign _0200_ = in_data[278] & _0025_;
  assign out_data[416] = _0272_ & _0604_;
  assign _0605_ = _0606_ & _0146_;
  assign _0032_ = _0122_ & _0084_;
  assign _0607_ = _0608_ & _0477_;
  assign _0549_ = _0610_ & _0609_;
  assign _0611_ = _0146_ & _0194_;
  assign _0612_ = _0594_ & _0270_;
  assign _0613_ = _0614_ & _0226_;
  assign _0157_ = _0153_ & _0015_;
  assign _0091_ = _0616_ & _0615_;
  assign _0198_ = _0065_ & _0617_;
  assign _0283_ = _0618_ & _0219_;
  assign _0619_ = _0241_ & _0620_;
  assign _0621_ = _0622_ & _0221_;
  assign _0246_ = _0320_ & _0108_;
  assign _0623_ = _0624_ & _0043_;
  assign _0180_ = _0625_ & _0251_;
  assign _0171_ = _0626_ & _0270_;
  assign _0627_ = _0628_ & _0175_;
  assign _0629_ = _0572_ & _0630_;
  assign _0631_ = _0057_ & _0401_;
  assign _0632_ = _0490_ & _0633_;
  assign _0101_ = _0025_ & in_data[679];
  assign _0634_ = _0228_ & _0055_;
  assign _0481_ = _0198_ & _0069_;
  assign _0455_ = _0071_ & _0241_;
  assign _0215_ = _0267_ & _0357_;
  assign _0635_ = _0636_ & _0412_;
  assign _0637_ = _0639_ & _0638_;
  assign _0640_ = _0138_ & _0082_;
  assign _0641_ = _0318_ & _0419_;
  assign _0552_ = _0143_ & _0642_;
  assign _0643_ = _0645_ & _0644_;
  assign _0646_ = _0647_ & _0419_;
  assign _0648_ = _0623_ & _0649_;
  assign _0650_ = _0625_ & _0651_;
  assign _0652_ = _0653_ & _0311_;
  assign _0654_ = _0572_ & _0112_;
  assign _0655_ = _0609_ & _0656_;
  assign _0657_ = _0401_ & _0565_;
  assign _0510_ = _0658_ & _0180_;
  assign _0659_ = _0609_ & _0565_;
  assign _0660_ = _0661_ & _0259_;
  assign _0662_ = _0248_ & _0469_;
  assign _0356_ = _0025_ & _0154_;
  assign _0663_ = _0309_ & _0453_;
  assign _0664_ = _0665_ & _0488_;
  assign _0666_ = _0668_ & _0667_;
  assign _0669_ = _0631_ & _0134_;
  assign _0071_ = _0197_ & _0152_;
  assign _0670_ = _0617_ & _0192_;
  assign _0296_ = _0316_ & _0671_;
  assign _0672_ = _0674_ & _0673_;
  assign _0675_ = _0677_ & _0676_;
  assign _0351_ = _0679_ & _0678_;
  assign _0680_ = _0615_ & _0620_;
  assign _0681_ = _0524_ & _0682_;
  assign _0307_ = _0684_ & _0683_;
  assign _0685_ = _0076_ & _0519_;
  assign _0686_ = _0572_ & _0687_;
  assign _0689_ = _0691_ & _0690_;
  assign _0484_ = _0140_ & _0692_;
  assign _0323_ = _0071_ & _0082_;
  assign _0694_ = _0225_ & _0661_;
  assign _0695_ = _0025_ & _0696_;
  assign _0525_ = _0697_ & _0228_;
  assign _0097_ = _0197_ & _0237_;
  assign _0456_ = _0071_ & _0363_;
  assign _0698_ = _0212_ & _0335_;
  assign _0699_ = _0700_ & _0069_;
  assign _0701_ = _0214_ & _0642_;
  assign _0406_ = _0702_ & _0332_;
  assign _0704_ = _0706_ & _0705_;
  assign _0707_ = _0709_ & _0708_;
  assign _0710_ = _0712_ & _0711_;
  assign _0464_ = _0134_ & _0272_;
  assign _0713_ = _0296_ & _0343_;
  assign _0714_ = _0563_ & _0217_;
  assign _0027_ = _0716_ & _0715_;
  assign _0717_ = _0167_ & _0662_;
  assign _0718_ = _0720_ & _0719_;
  assign _0721_ = _0401_ & _0722_;
  assign _0723_ = _0595_ & _0165_;
  assign out_data[1184] = _0725_ & _0724_;
  assign _0727_ = _0102_ & _0728_;
  assign _0729_ = _0730_ & _0565_;
  assign _0731_ = _0733_ & _0732_;
  assign _0636_ = _0529_ & _0734_;
  assign _0735_ = _0321_ & _0736_;
  assign _0019_ = _0737_ & _0071_;
  assign _0738_ = _0739_ & _0641_;
  assign _0741_ = _0034_ & _0239_;
  assign _0743_ = _0744_ & _0590_;
  assign _0745_ = _0746_ & _0148_;
  assign _0747_ = _0148_ & _0295_;
  assign _0088_ = _0018_ & _0748_;
  assign _0749_ = _0613_ & _0750_;
  assign _0751_ = _0752_ & _0248_;
  assign _0753_ = _0241_ & _0134_;
  assign _0754_ = _0756_ & _0755_;
  assign _0757_ = _0689_ & _0758_;
  assign _0518_ = _0033_ & _0287_;
  assign _0761_ = _0717_ & _0762_;
  assign _0763_ = _0765_ & _0764_;
  assign _0768_ = _0038_ & _0454_;
  assign _0770_ = _0771_ & _0152_;
  assign _0769_ = _0317_ & _0226_;
  assign _0772_ = _0663_ & _0773_;
  assign _0203_ = _0221_ & _0277_;
  assign _0774_ = _0598_ & _0775_;
  assign _0776_ = _0778_ & _0777_;
  assign _0780_ = _0782_ & _0781_;
  assign _0783_ = _0784_ & _0145_;
  assign _0354_ = _0529_ & _0690_;
  assign _0786_ = _0663_ & _0787_;
  assign _0788_ = _0619_ & _0789_;
  assign _0079_ = _0792_ & _0784_;
  assign _0796_ = _0379_ & _0736_;
  assign _0159_ = _0025_ & _0359_;
  assign _0797_ = _0799_ & _0798_;
  assign _0800_ = _0801_ & _0387_;
  assign _0379_ = _0150_ & _0317_;
  assign _0802_ = _0094_ & _0803_;
  assign _0804_ = _0806_ & _0805_;
  assign _0807_ = _0808_ & _0317_;
  assign _0085_ = _0111_ & _0295_;
  assign _0809_ = _0212_ & _0453_;
  assign _0810_ = _0812_ & _0811_;
  assign _0813_ = _0640_ & _0735_;
  assign _0814_ = _0743_ & _0408_;
  assign _0815_ = _0816_ & _0134_;
  assign _0820_ = _0373_ & _0797_;
  assign _0821_ = _0113_ & _0221_;
  assign _0823_ = _0776_ & _0328_;
  assign _0824_ = _0826_ & _0825_;
  assign _0827_ = _0046_ & _0828_;
  assign _0446_ = _0450_ & _0829_;
  assign _0210_ = _0633_ & _0316_;
  assign _0831_ = _0833_ & _0832_;
  assign _0834_ = _0392_ & _0835_;
  assign _0837_ = _0838_ & _0309_;
  assign _0843_ = _0845_ & _0844_;
  assign _0846_ = _0848_ & _0847_;
  assign _0527_ = _0274_ & _0852_;
  assign _0856_ = _0636_ & _0857_;
  assign _0858_ = _0860_ & _0859_;
  assign _0861_ = _0863_ & _0862_;
  assign _0867_ = _0869_ & _0868_;
  assign _0870_ = _0757_ & _0178_;
  assign _0573_ = _0189_ & _0864_;
  assign _0522_ = _0609_ & _0069_;
  assign _0876_ = _0878_ & _0877_;
  assign _0884_ = _0885_ & _0640_;
  assign _0886_ = _0888_ & _0887_;
  assign _0902_ = _0904_ & _0903_;
  assign _0905_ = _0908_ & _0907_;
  assign _0911_ = ~((_0890_ & _0912_) | _0209_);
  assign _0917_ = ~((_0639_ & _0582_) | _0600_);
  assign _0502_ = ~((_0918_ & _0359_) | _0033_);
  assign _0919_ = ~((_0111_ & _0920_) | _0033_);
  assign _0543_ = ~((_0258_ & _0922_) | _0921_);
  assign _0049_ = ~((_0926_ & _0925_) | _0228_);
  assign _0931_ = ~((_0698_ & _0018_) | _0273_);
  assign _0933_ = ~((_0935_ & _0271_) | _0934_);
  assign _0599_ = ~((_0325_ & _0748_) | _0752_);
  assign _0228_ = ~((_0096_ & _0238_) | _0096_);
  assign _0950_ = ~((_0953_ & _0952_) | _0951_);
  assign _0955_ = ~((_0957_ & _0956_) | _0675_);
  assign _0959_ = ~((_0962_ & _0961_) | _0960_);
  assign _0964_ = ~((_0837_ & _0812_) | _0965_);
  assign out_data[1312] = ~((_0977_ & _0110_) | _0009_);
  assign out_data[960] = ~((_0111_ & _0856_) | _0069_);
  assign out_data[864] = ~((_0980_ & _0979_) | _0978_);
  assign out_data[768] = ~((_0982_ & _0034_) | _0981_);
  assign _0873_ = ~((_0039_ & _0434_) | _0022_);
  assign _0046_ = ~((_0019_ & _0661_) | _0983_);
  assign _0984_ = ~((_0205_ & _0985_) | _0159_);
  assign _0289_ = ~((_0067_ & _0113_) | _0986_);
  assign _0357_ = ~((_0690_ & _0136_) | _0065_);
  assign _0987_ = ~((_0586_ & _0988_) | _0141_);
  assign _0082_ = ~((_0154_ & _0033_) | _0152_);
  assign _0208_ = ~((_0101_ & _0775_) | _0599_);
  assign _0278_ = ~((_0989_ & _0318_) | _0419_);
  assign _0178_ = ~((_0277_ & _0096_) | _0490_);
  assign _0811_ = ~((_0101_ & _0058_) | _0191_);
  assign _0665_ = ~((_0043_ & _0206_) | _0990_);
  assign _0991_ = ~((_0994_ & _0993_) | _0992_);
  assign _0316_ = ~((_0103_ & _0993_) | _0529_);
  assign _0454_ = ~((_0383_ & _0137_) | _0206_);
  assign _0995_ = ~((_0636_ & _0317_) | _0611_);
  assign _0841_ = ~((_0065_ & _0626_) | _0098_);
  assign _0249_ = ~((_0962_ & _0000_) | _0996_);
  assign _0212_ = ~((_0055_ & _0615_) | _0210_);
  assign _0997_ = ~((_0999_ & _0316_) | _0998_);
  assign _0412_ = ~((_0058_ & _0164_) | _1000_);
  assign _1001_ = ~((_0258_ & _0109_) | _1002_);
  assign _1003_ = ~((_0891_ & _0289_) | _0235_);
  assign _1004_ = ~((_0065_ & _0594_) | _0136_);
  assign _1005_ = ~((_0113_ & _0228_) | _0104_);
  assign _0915_ = ~((_0149_ & _0356_) | _0022_);
  assign _0035_ = ~((_0194_ & _0151_) | _0095_);
  assign _1006_ = ~((_0152_ & _1007_) | _0485_);
  assign _0785_ = ~((_0175_ & _0177_) | _0591_);
  assign _0425_ = ~((_0166_ & _0250_) | _1008_);
  assign _0808_ = ~((_0637_ & _1010_) | _1009_);
  assign _0503_ = ~((_0801_ & _1012_) | _1011_);
  assign _0793_ = ~((_0589_ & _0117_) | _0012_);
  assign _1013_ = ~((_0611_ & _0989_) | _1014_);
  assign _1015_ = ~((_0175_ & _0988_) | _1016_);
  assign _0214_ = ~((_1017_ & _0354_) | _0620_);
  assign _0683_ = ~((_0139_ & _0213_) | _0609_);
  assign _1018_ = ~((_0140_ & _0242_) | _0251_);
  assign _1019_ = ~((_0919_ & _0343_) | _0272_);
  assign _1020_ = ~((_0019_ & _0537_) | _0121_);
  assign out_data[1920] = ~((_0645_ & _1021_) | _0116_);
  assign _0340_ = ~((_0149_ & _0529_) | _1022_);
  assign _1023_ = ~((_0057_ & _1024_) | _0678_);
  assign _0376_ = ~((_0671_ & _0755_) | _0272_);
  assign _0369_ = ~((_0251_ & _0065_) | _0227_);
  assign _1025_ = ~((_0615_ & _1014_) | _1026_);
  assign out_data[1344] = ~((_1028_ & _0097_) | _1027_);
  assign _0865_ = ~((_1030_ & _1029_) | _0936_);
  assign _1031_ = ~((_0003_ & _0094_) | _1032_);
  assign _1033_ = ~((_0625_ & _0108_) | _0091_);
  assign _0914_ = ~((_0304_ & _1020_) | _0979_);
  assign _0322_ = ~((_1034_ & _0613_) | _0469_);
  assign _1035_ = ~((_0202_ & out_data[1344]) | _0316_);
  assign _1036_ = ~((_0264_ & _0458_) | _1037_);
  assign _1038_ = ~((_1039_ & _0171_) | _0590_);
  assign _0732_ = ~((_1041_ & _0151_) | _1040_);
  assign _0682_ = ~((_0283_ & _0692_) | _0211_);
  assign _0475_ = ~((_0255_ & _0655_) | _0623_);
  assign _0311_ = ~((_1042_ & _0043_) | _0918_);
  assign _1043_ = ~((_0187_ & _1044_) | _0015_);
  assign _0687_ = ~((_0873_ & _0264_) | _1045_);
  assign _0835_ = ~((_0096_ & _0042_) | _0481_);
  assign _0191_ = ~((_0103_ & _1046_) | _0311_);
  assign _0463_ = ~((_0306_ & _0134_) | _1046_);
  assign _1047_ = ~((_0117_ & _0143_) | _0529_);
  assign _0532_ = ~((_0984_ & _0700_) | _1048_);
  assign _1051_ = ~((_0454_ & _0199_) | _0044_);
  assign _1052_ = ~((_0726_ & _0612_) | _0671_);
  assign _1053_ = ~((_0615_ & _0389_) | _1054_);
  assign _1055_ = ~((_0219_ & _1056_) | _0525_);
  assign _0890_ = ~((_0043_ & _0675_) | _0082_);
  assign _1057_ = ~((_0219_ & _0593_) | _1058_);
  assign _1061_ = ~((_1020_ & _0161_) | _1062_);
  assign _1063_ = ~((_0016_ & _0096_) | _0593_);
  assign _1065_ = ~((_0292_ & _1066_) | _0924_);
  assign _1067_ = ~((_1069_ & _0726_) | _1068_);
  assign _1073_ = ~((_0525_ & _0454_) | _1074_);
  assign _1075_ = ~((_1061_ & _0922_) | _0713_);
  assign _0058_ = ~((_0318_ & _0733_) | _0084_);
  assign _1076_ = ~((_1078_ & _1077_) | _0631_);
  assign _0562_ = ~((_0128_ & _1082_) | _1081_);
  assign _0897_ = ~((_1083_ & _1061_) | _0489_);
  assign _1084_ = ~((_0134_ & _0134_) | _0003_);
  assign _1085_ = ~((_1087_ & _1086_) | _0752_);
  assign _1088_ = ~((_0941_ & _0123_) | _0205_);
  assign _1089_ = ~((_0901_ & _1090_) | _0000_);
  assign _0756_ = ~((_0692_ & _0490_) | _1091_);
  assign _1092_ = ~((_1093_ & _0312_) | _0856_);
  assign _1095_ = ~((_0692_ & _1097_) | _1096_);
  assign _1098_ = ~((_1100_ & _0578_) | _1099_);
  assign _0116_ = ~((_0343_ & _0610_) | _0096_);
  assign _0838_ = ~((_1101_ & _0353_) | _0161_);
  assign _1102_ = ~((_1104_ & _1103_) | _0505_);
  assign _0609_ = ~((_0265_ & _0311_) | _0238_);
  assign _1105_ = ~((_1107_ & _1106_) | _0419_);
  assign _1108_ = ~((_0134_ & _1109_) | _0795_);
  assign _1110_ = ~((_0915_ & _1056_) | _1111_);
  assign _0875_ = ~((_0662_ & _1056_) | _0134_);
  assign _1112_ = ~((_0335_ & _1113_) | _0166_);
  assign _0805_ = ~((_0057_ & _0708_) | _0531_);
  assign _0497_ = ~((_0170_ & _1115_) | _0740_);
  assign _0083_ = ~((_0503_ & _0565_) | _0434_);
  assign _0416_ = ~((_0278_ & _0164_) | _0269_);
  assign _1116_ = ~((_0617_ & _0727_) | _0787_);
  assign _0371_ = ~((_0891_ & _1119_) | _0259_);
  assign _1120_ = ~((_0152_ & _0370_) | _0145_);
  assign _0752_ = ~((_0237_ & _0116_) | _0232_);
  assign _0829_ = ~((_0825_ & _0854_) | _0270_);
  assign _1123_ = ~((_0731_ & _1124_) | _0598_);
  assign _1125_ = ~((_0572_ & _1117_) | _1126_);
  assign _0146_ = ~((_0609_ & _0306_) | _0464_);
  assign _0913_ = ~((_1127_ & _0157_) | _0733_);
  assign _0859_ = ~((_1131_ & _1130_) | _0866_);
  assign _1133_ = ~((_0774_ & _1110_) | _0348_);
  assign _1135_ = ~((_1137_ & out_data[1344]) | _1136_);
  assign _1139_ = ~((_1141_ & _1140_) | _0697_);
  assign _1142_ = ~((_1143_ & _1013_) | _0854_);
  assign _0422_ = ~((_1146_ & _0838_) | _1145_);
  assign _0860_ = ~((_0455_ & _0726_) | _1147_);
  assign _1148_ = ~((_0109_ & _1072_) | _0166_);
  assign _1149_ = ~((_0071_ & _0228_) | _1150_);
  assign _1151_ = ~((_1153_ & _0101_) | _1152_);
  assign _1154_ = ~((_0871_ & _1156_) | _1155_);
  assign _0478_ = ~((_1158_ & _0217_) | _1157_);
  assign _0430_ = ~((_0341_ & _0044_) | _0578_);
  assign _1165_ = ~((_0631_ & _1166_) | _0102_);
  assign _0603_ = ~((_0294_ & _0401_) | _0134_);
  assign _1169_ = ~((_1170_ & _1025_) | _0096_);
  assign _1170_ = ~((_0290_ & _0586_) | _0733_);
  assign _0555_ = ~((_0821_ & _1174_) | _1173_);
  assign _1177_ = ~((_0249_ & _0343_) | _0443_);
  assign _0957_ = ~((_1180_ & _0860_) | _0947_);
  assign _1181_ = ~((_0569_ & _1182_) | _0841_);
  assign _1183_ = ~((_1170_ & _1184_) | _0062_);
  assign _0361_ = ~((_0316_ & _0152_) | _0490_);
  assign _1186_ = ~((_1187_ & _0355_) | _0109_);
  assign _1188_ = ~((_0014_ & _0994_) | _0212_);
  assign _1190_ = ~((_0605_ & _0361_) | _0096_);
  assign _0507_ = ~((_0770_ & _1192_) | _1191_);
  assign _1196_ = ~((_0958_ & _1025_) | _1036_);
  assign _0934_ = ~((_1200_ & _1199_) | _1198_);
  assign _0581_ = ~((_0152_ & _1202_) | _1201_);
  assign _1205_ = ~((_0096_ & _0304_) | _1206_);
  assign _1207_ = ~((_1208_ & _1177_) | _1005_);
  assign _0617_ = ~((_1211_ & _0625_) | _1210_);
  assign _1212_ = ~((_0261_ & _1213_) | _0058_);
  assign _1215_ = ~((_0867_ & _1217_) | _1216_);
  assign _1218_ = ~((_0245_ & _0885_) | _0038_);
  assign _0975_ = ~((_1219_ & _0337_) | _0932_);
  assign _1220_ = ~((_1222_ & _0898_) | _1221_);
  assign _0960_ = ~((_1223_ & _0502_) | _0993_);
  assign _1229_ = ~((_0400_ & _0689_) | _1230_);
  assign _1234_ = ~((_0671_ & _1235_) | _1199_);
  assign _1237_ = ~((_1241_ & _1240_) | (_1239_ & _1238_));
  assign _0090_ = ~((_0600_ & _0670_) | (_0539_ & _1246_));
  assign _0059_ = ~((_1255_ & _0149_) | (_0606_ & _1253_));
  assign _1259_ = ~((_0649_ & _1028_) | (_0305_ & _0389_));
  assign _0434_ = ~((_0116_ & _1016_) | (_0529_ & _0887_));
  assign _1264_ = ~((_0672_ & _0191_) | (_0110_ & _1265_));
  assign _1266_ = ~((_1170_ & _0250_) | (_0039_ & _0134_));
  assign _1275_ = ~((_1188_ & _0505_) | (_0286_ & _0099_));
  assign _0057_ = ~((_0071_ & _0306_) | (_1278_ & _1276_));
  assign _0094_ = ~((_1284_ & _1283_) | (_0097_ & _1282_));
  assign _1289_ = ~((_0195_ & _0183_) | (_1290_ & _0546_));
  assign _0591_ = ~((_0044_ & _0463_) | (_0200_ & _0625_));
  assign _0982_ = ~((_0582_ & _0861_) | (_0248_ & _0732_));
  assign out_data[1856] = ~((_0554_ & _1028_) | (_1265_ & _1292_));
  assign out_data[1824] = ~((_1294_ & _0295_) | (_0416_ & _1293_));
  assign out_data[1792] = ~((_1265_ & _1297_) | (_1296_ & _1295_));
  assign out_data[1760] = ~((_0830_ & _0931_) | (_1298_ & _0406_));
  assign out_data[1728] = ~((_0080_ & _0879_) | (_0565_ & _1209_));
  assign out_data[1696] = ~((_1300_ & _0457_) | (_1299_ & _0639_));
  assign out_data[1632] = ~((_0051_ & _1301_) | (_0480_ & _1212_));
  assign _1302_ = ~((_0325_ & _0265_) | (_0044_ & _0272_));
  assign out_data[736] = ~((_0834_ & _1303_) | (_0420_ & _0636_));
  assign out_data[160] = ~((_0134_ & out_data[64]) | (_0057_ & _1304_));
  assign _0801_ = ~((_1306_ & _0203_) | (_0191_ & _1305_));
  assign _0469_ = ~((_1307_ & _1000_) | (_0468_ & _1046_));
  assign _1113_ = ~((_1310_ & _1309_) | (_1308_ & _0197_));
  assign _1311_ = ~((_0438_ & _0905_) | (_1312_ & _0121_));
  assign _0359_ = ~((_1000_ & _0101_) | (_0033_ & _1000_));
  assign _0163_ = ~((_1313_ & _0581_) | (_0096_ & _0125_));
  assign _0139_ = ~((_0177_ & _0752_) | (_1314_ & _0563_));
  assign _1315_ = ~((_0094_ & _1113_) | (_0121_ & _0219_));
  assign _0055_ = ~((_0272_ & _1316_) | (_0318_ & _0149_));
  assign _0989_ = ~((_1318_ & _0099_) | (_0600_ & _1317_));
  assign _1027_ = ~((_0529_ & _0206_) | (_0524_ & _0097_));
  assign _0332_ = ~((_0469_ & _0343_) | (_1320_ & _1319_));
  assign _0651_ = ~((_1321_ & _0602_) | (_0317_ & _0419_));
  assign _0489_ = ~((_0043_ & _0605_) | (_0175_ & _0058_));
  assign _1322_ = ~((_1323_ & _0065_) | (_0661_ & _1000_));
  assign _0909_ = ~((_0615_ & _1326_) | (_1325_ & _1324_));
  assign _0348_ = ~((_1206_ & _0651_) | (_0994_ & _1283_));
  assign _0540_ = ~((_0915_ & _0019_) | (_0289_ & _0259_));
  assign _0231_ = ~((_0016_ & _0612_) | (_0801_ & _0325_));
  assign _1127_ = ~((_1327_ & _0019_) | (_0335_ & _0205_));
  assign _0401_ = ~((_0103_ & _1328_) | (_0228_ & _0513_));
  assign _1329_ = ~((_0139_ & _0071_) | (_1330_ & _0212_));
  assign _0242_ = ~((_0250_ & _0221_) | (_0281_ & _0613_));
  assign _0306_ = ~((_0128_ & _0403_) | (_0043_ & _0150_));
  assign _1028_ = ~((_0152_ & _0134_) | (_0489_ & _0529_));
  assign _1331_ = ~((_0152_ & _0231_) | (_1332_ & _0043_));
  assign _0186_ = ~((_0009_ & _0025_) | (_0129_ & _1333_));
  assign _0733_ = ~((in_data[103] & _0317_) | (_0149_ & _0127_));
  assign _1334_ = ~((_1335_ & _0219_) | (_0116_ & _0135_));
  assign _1336_ = ~((_1338_ & _0133_) | (_0529_ & _1337_));
  assign _0411_ = ~((_0000_ & _0144_) | (_0623_ & _0733_));
  assign _0816_ = ~((_1003_ & _1334_) | (_0454_ & _0989_));
  assign _1339_ = ~((_0168_ & _0204_) | (_1027_ & _0023_));
  assign _0076_ = ~((_0199_ & _0112_) | (_1340_ & _0095_));
  assign _1056_ = ~((_1341_ & _0502_) | (_0716_ & _0067_));
  assign _1342_ = ~((_0899_ & _1344_) | (_0420_ & _1343_));
  assign _1345_ = ~((_0979_ & _0053_) | (_0918_ & _0299_));
  assign _1017_ = ~((_0611_ & _0166_) | (_0080_ & _1334_));
  assign _1347_ = ~((_1350_ & _1349_) | (_1348_ & _0401_));
  assign _0789_ = ~((_0164_ & _0309_) | (_0042_ & _0489_));
  assign _1046_ = ~((_1351_ & _0189_) | (_0134_ & _1346_));
  assign _0385_ = ~((_0303_ & _1352_) | (_0170_ & _0692_));
  assign _0460_ = ~((_1001_ & _0438_) | (_0272_ & _0598_));
  assign _1021_ = ~((_1354_ & _1353_) | (_0080_ & _0134_));
  assign _0490_ = ~((_1355_ & _0101_) | (_0101_ & _0125_));
  assign _1024_ = ~((_0110_ & _0019_) | (_0317_ & _1026_));
  assign _1356_ = ~((_0999_ & _0175_) | (_1357_ & _0032_));
  assign _0386_ = ~((_0018_ & _0081_) | (_0401_ & _0082_));
  assign _0237_ = ~((_0915_ & _0529_) | (_0915_ & _0573_));
  assign _1358_ = ~((_0207_ & _0489_) | (_1360_ & _1359_));
  assign _0394_ = ~((_0620_ & _1362_) | (_1361_ & _0113_));
  assign _0084_ = ~((_0359_ & _0043_) | (_0200_ & _0232_));
  assign _1363_ = ~((_0082_ & _1086_) | (_1364_ & _0984_));
  assign _1096_ = ~((_0454_ & _1365_) | (_1225_ & _0229_));
  assign _1366_ = ~((_0289_ & _0094_) | (_1367_ & _0566_));
  assign _0197_ = ~((_0134_ & _0529_) | (_0241_ & _0205_));
  assign _1114_ = ~((_0613_ & _0613_) | (_1368_ & _0065_));
  assign _0794_ = ~((_0105_ & _1336_) | (_0997_ & _1131_));
  assign _0830_ = ~((_0274_ & _0190_) | (_1369_ & _0350_));
  assign _1370_ = ~((_1001_ & _0146_) | (_0316_ & _0411_));
  assign _1371_ = ~((_0626_ & _0246_) | (_0672_ & _1372_));
  assign _0269_ = ~((_0848_ & _0690_) | (_0489_ & _0196_));
  assign _1161_ = ~((_1147_ & _0635_) | (_0231_ & _1373_));
  assign _0759_ = ~((_0841_ & _0726_) | (_1374_ & _0238_));
  assign _0417_ = ~((_0112_ & _1136_) | (_0193_ & _0490_));
  assign _1375_ = ~((_0748_ & _1376_) | (_1331_ & _1360_));
  assign _1377_ = ~((_0656_ & _0619_) | (_1379_ & _1378_));
  assign _1380_ = ~((_1382_ & _0133_) | (_1381_ & _1056_));
  assign _1283_ = ~((_1384_ & _0127_) | (_0275_ & _1383_));
  assign _0285_ = ~((_0726_ & _0206_) | (_0519_ & _0134_));
  assign _0904_ = ~((_0243_ & _1387_) | (_1386_ & _1385_));
  assign _1388_ = ~((_1389_ & _0488_) | (_0984_ & _0523_));
  assign _1390_ = ~((_0263_ & _0946_) | (_0201_ & _1391_));
  assign _0138_ = ~((_1034_ & _0033_) | (_0915_ & _0152_));
  assign _1392_ = ~((_0629_ & _0586_) | (_0096_ & _1393_));
  assign _1394_ = ~((_0217_ & _0014_) | (_0238_ & _0919_));
  assign _1395_ = ~((_1397_ & _1396_) | (_1077_ & _0161_));
  assign _0338_ = ~((_0191_ & _1381_) | (_0096_ & _0062_));
  assign _0941_ = ~((_0794_ & _0217_) | (_1398_ & _0565_));
  assign _0901_ = ~((_0502_ & _0622_) | (_0221_ & _1375_));
  assign _1399_ = ~((_1017_ & _0795_) | (_0678_ & _0149_));
  assign _0586_ = ~((_0529_ & _0194_) | (_0237_ & _0043_));
  assign _1208_ = ~((_1400_ & _0502_) | (_0254_ & _1302_));
  assign _0524_ = ~((_0529_ & in_data[928]) | (_0316_ & in_data[2096]));
  assign _1401_ = ~((_0149_ & _1403_) | (_0306_ & _1402_));
  assign _0894_ = ~((_0402_ & _1404_) | (_0065_ & _0450_));
  assign _0799_ = ~((_1407_ & _0711_) | (_1406_ & _1405_));
  assign _0784_ = ~((_0255_ & _0995_) | (_0239_ & _1028_));
  assign _0270_ = ~((_0033_ & _0134_) | (_0993_ & _0018_));
  assign _0467_ = ~((_0013_ & _0214_) | (_1034_ & _1072_));
  assign _0888_ = ~((_1408_ & _0936_) | (_0222_ & _0403_));
  assign _1409_ = ~((_0316_ & _1410_) | (_1147_ & _0455_));
  assign _0866_ = ~((_0258_ & _1342_) | (_0043_ & _0368_));
  assign _1411_ = ~((_0258_ & _0128_) | (_0288_ & _1412_));
  assign _0977_ = ~((_0337_ & _0905_) | (_0759_ & _0307_));
  assign _0560_ = ~((_0091_ & _0065_) | (_0505_ & _0109_));
  assign _0740_ = ~((_1413_ & _0080_) | (_0039_ & _1245_));
  assign _0766_ = ~((_0627_ & _0044_) | (_0572_ & _0419_));
  assign _0530_ = ~((_0879_ & _1417_) | (_0065_ & _0385_));
  assign _1418_ = ~((_0097_ & _0799_) | (_0335_ & _0175_));
  assign _0758_ = ~((_1419_ & _0190_) | (_0012_ & _0578_));
  assign _0342_ = ~((_0052_ & _1339_) | (_0247_ & _1420_));
  assign _1393_ = ~((_0106_ & _0403_) | (_0401_ & _0101_));
  assign _1422_ = ~((_0594_ & _1423_) | (_0160_ & _0263_));
  assign _1424_ = ~((_0368_ & _0057_) | (_0032_ & _0726_));
  assign _1301_ = ~((_1426_ & _0708_) | (_0641_ & _0242_));
  assign _0433_ = ~((_1428_ & _0385_) | (_1427_ & _1028_));
  assign _0353_ = ~((_1430_ & _1406_) | (_1429_ & _0289_));
  assign _0907_ = ~((_0318_ & _0228_) | (_0610_ & _0317_));
  assign _1433_ = ~((_0150_ & _0351_) | (_1170_ & _1406_));
  assign _1434_ = ~((_0287_ & _1147_) | (_1053_ & _0450_));
  assign _1435_ = ~((_0193_ & _0337_) | (_0191_ & _1056_));
  assign _0608_ = ~((_0082_ & _0022_) | (_0993_ & _0152_));
  assign _1438_ = ~((_1347_ & _0159_) | (_0175_ & _1147_));
  assign _1439_ = ~((_1345_ & _0287_) | (_0729_ & _1440_));
  assign _1224_ = ~((_1442_ & _0755_) | (_0537_ & _0890_));
  assign _1443_ = ~((_1053_ & _1434_) | (_1444_ & _1409_));
  assign _1290_ = ~((_1379_ & _1446_) | (_1445_ & _1164_));
  assign _0064_ = ~((_1448_ & _1447_) | (_0235_ & _1056_));
  assign _1137_ = ~((_0537_ & _0590_) | (_0292_ & _1076_));
  assign _1451_ = ~((_0436_ & _0202_) | (_1452_ & _0179_));
  assign _0033_ = ~((_0241_ & _0200_) | (_0025_ & _0356_));
  assign _1454_ = ~((_0434_ & _0953_) | (_1456_ & _1455_));
  assign _1457_ = ~((_1436_ & _0190_) | (_1458_ & _0116_));
  assign _1459_ = ~((_0825_ & _1290_) | (_1460_ & _0194_));
  assign _1462_ = ~((_0192_ & _0915_) | (_0146_ & _0599_));
  assign _1299_ = ~((_0144_ & _0924_) | (_0615_ & _0096_));
  assign _1463_ = ~((_0717_ & _1464_) | (_0134_ & _0009_));
  assign _1465_ = ~((_0299_ & _0046_) | (_1466_ & _1384_));
  assign _1471_ = ~((_1472_ & _0032_) | (_0243_ & _1187_));
  assign _1473_ = ~((_1047_ & _0949_) | (_1474_ & _1395_));
  assign _0050_ = ~((_1477_ & _0855_) | (_1025_ & _1017_));
  assign _1478_ = ~((_1480_ & _1004_) | (_0784_ & _1479_));
  assign _1481_ = ~((_0615_ & _0469_) | (_1000_ & _1019_));
  assign _1228_ = ~((_0082_ & _0907_) | (_0091_ & _0175_));
  assign _0103_ = ~((_0104_ & _1476_) | (_1467_ & _0189_));
  assign _1129_ = ~((_0637_ & _0117_) | (_1089_ & _0589_));
  assign _1486_ = ~((_1488_ & _1487_) | (_0279_ & _0490_));
  assign _1491_ = ~((_1493_ & _1492_) | (_0656_ & _0699_));
  assign _1497_ = ~((_0712_ & _0394_) | (_0718_ & _0548_));
  assign _1178_ = ~((_0187_ & _1500_) | (_0097_ & _0778_));
  assign _1197_ = ~((_0134_ & _0785_) | (_1066_ & _0697_));
  assign _1501_ = ~((_0672_ & _1502_) | (_0115_ & _0800_));
  assign _1362_ = ~((_0058_ & _0082_) | (_0383_ & _0402_));
  assign out_data[256] = ~((_1197_ & _0694_) | (_1505_ & _0228_));
  assign _0639_ = ~((_0320_ & _0132_) | (_0228_ & _1507_));
  assign _0571_ = ~((_0548_ & _0119_) | (_0050_ & _1509_));
  assign _0193_ = ~((_0068_ & _1283_) | (_0356_ & _0219_));
  assign _0443_ = ~((_0218_ & _0690_) | (_0019_ & _0245_));
  assign _0739_ = ~((_0106_ & _0733_) | (_0127_ & _0127_));
  assign _1512_ = ~((_0753_ & _0738_) | (_0989_ & _1513_));
  assign _0039_ = ~((_0463_ & _0287_) | (_1511_ & _0383_));
  assign _1514_ = ~((_1515_ & _0137_) | (_0461_ & _1224_));
  assign _0885_ = ~((_0620_ & _0042_) | (_1517_ & _1516_));
  assign _1158_ = ~((_0012_ & _1519_) | (_0237_ & _0811_));
  assign _0857_ = ~((_1521_ & _1520_) | (_0690_ & _0128_));
  assign _0575_ = ~((_1524_ & _1171_) | (_1523_ & _1522_));
  assign _1527_ = ~((_0769_ & _0152_) | (_0356_ & _0250_));
  assign _0486_ = ~((_0134_ & _1529_) | (_0725_ & _0856_));
  assign _0947_ = ~((_0412_ & _0317_) | (_1533_ & _1532_));
  assign _0044_ = ~((_0227_ & _0639_) | (_0315_ & _0609_));
  assign _0963_ = ~((_1053_ & _1539_) | (_1538_ & _1537_));
  assign _1257_ = ~((_1545_ & _1544_) | (_0490_ & _1543_));
  assign _0001_ = ~((_0228_ & _1547_) | (_0914_ & _1368_));
  assign _0144_ = ~((_1362_ & _0304_) | (_0193_ & _0311_));
  assign _0043_ = ~((_0356_ & _0356_) | (_0319_ & _0127_));
  assign _1555_ = ~((_1556_ & _0527_) | (_0176_ & _0282_));
  assign _1557_ = ~((_0325_ & _0905_) | (_0799_ & _1558_));
  assign _0961_ = ~((_0435_ & _1299_) | (_0257_ & _0944_));
  assign _0515_ = ~((_1148_ & _1057_) | (_0071_ & _1561_));
  assign _0582_ = ~((_0772_ & _1571_) | (_1570_ & _0431_));
  assign _0565_ = ~((_0408_ & _1569_) | (_1568_ & _0150_));
  assign _1239_ = ~((_0559_ & _1183_) | (_1573_ & _0201_));
  assign _1574_ = ~((_1196_ & _0900_) | (_1501_ & _1575_));
  assign _0534_ = ~((_1584_ & _0831_) | (_0726_ & _1583_));
  assign _1587_ = ~((_1588_ & _1199_) | (_0816_ & _0787_));
  assign _1589_ = ~((_0134_ & _0907_) | (_0272_ & _1590_));
  assign _0887_ = ~((_0111_ & _0464_) | (_1309_ & _1136_));
  assign _1599_ = ~((_0816_ & _1557_) | (_1600_ & _0745_));
  assign _0951_ = ~((_1601_ & _1142_) | (_0148_ & _1137_));
  assign _0551_ = ~((_1603_ & _0437_) | (_0125_ & _1602_));
  assign _1648_ = _1649_ | _0486_;
  assign _1629_ = _0721_ | _1025_;
  assign _0226_ = _0356_ | _0238_;
  assign _1650_ = _1112_ | _1651_;
  assign _1657_ = _1607_ | _1658_;
  assign _1659_ = _1624_ | _0218_;
  assign _1660_ = _1399_ | _1661_;
  assign _0438_ = _0573_ | _0529_;
  assign _0678_ = _0130_ | _0359_;
  assign _1664_ = _0371_ | _0783_;
  assign _0936_ = _0146_ | _0084_;
  assign _0018_ = _0025_ | in_data[932];
  assign out_data[1216] = _0469_ | _0521_;
  assign out_data[576] = _0047_ | _0707_;
  assign _0013_ = _0306_ | _0893_;
  assign _0592_ = _0354_ | _0356_;
  assign _0781_ = _0521_ | _0356_;
  assign _0692_ = _1666_ | _0082_;
  assign _0477_ = _0642_ | _0025_;
  assign _0795_ = _0769_ | _0453_;
  assign _1130_ = _0193_ | _1315_;
  assign _0016_ = _0123_ | _0343_;
  assign _0700_ = _1211_ | _1136_;
  assign _0626_ = _0856_ | _0586_;
  assign _0848_ = _0205_ | _0046_;
  assign _1064_ = _1668_ | _1667_;
  assign _1247_ = _0625_ | _1669_;
  assign _0185_ = _0105_ | _0274_;
  assign _0267_ = _0324_ | _0716_;
  assign _1352_ = _0994_ | _0309_;
  assign _0000_ = _0645_ | _1393_;
  assign _0286_ = _1670_ | _0200_;
  assign _0854_ = _0152_ | _0988_;
  assign _0488_ = _1671_ | _0043_;
  assign _1449_ = _0325_ | _1322_;
  assign _0204_ = _1046_ | _0208_;
  assign _1391_ = _1672_ | _1483_;
  assign _0715_ = _0317_ | _0464_;
  assign _0034_ = _0152_ | _1069_;
  assign _1518_ = _0136_ | _0988_;
  assign _0436_ = _0328_ | _0848_;
  assign _0022_ = _0359_ | _0128_;
  assign _1134_ = _0025_ | _0265_;
  assign _0196_ = _0042_ | _0250_;
  assign _0730_ = _0656_ | _0055_;
  assign _0303_ = _0612_ | _0619_;
  assign _1144_ = _1005_ | _0032_;
  assign _1086_ = _1003_ | _1674_;
  assign _1245_ = _0228_ | _0175_;
  assign _0320_ = _0356_ | _1000_;
  assign _0448_ = _0106_ | _1673_;
  assign _0978_ = _0678_ | _0278_;
  assign _1663_ = _0690_ | _0317_;
  assign _1675_ = _0041_ | _0025_;
  assign _1235_ = _0152_ | _0022_;
  assign _0537_ = _0891_ | _0201_;
  assign _1026_ = _0135_ | _1518_;
  assign _1627_ = _0994_ | _0915_;
  assign _1066_ = _1676_ | _0250_;
  assign _0953_ = _0488_ | _0299_;
  assign _0671_ = _0438_ | _0042_;
  assign _0918_ = _0915_ | _0025_;
  assign _0638_ = _0025_ | _1677_;
  assign _0702_ = _0873_ | _0379_;
  assign _0505_ = _0769_ | _1678_;
  assign _0301_ = _1679_ | _0600_;
  assign _1680_ = _0193_ | _0454_;
  assign _1651_ = _0463_ | _0018_;
  assign _1425_ = _0203_ | _1681_;
  assign _0703_ = _0206_ | _1682_;
  assign _1174_ = _0654_ | _0116_;
  assign _1304_ = _0289_ | _1683_;
  assign _1128_ = _0250_ | _1684_;
  assign _0967_ = _0357_ | _0227_;
  assign _0724_ = _0148_ | _0703_;
  assign _0709_ = _0251_ | _0158_;
  assign _0221_ = _1255_ | _0915_;
  assign _0447_ = _0354_ | _1685_;
  assign _1686_ = _0436_ | _0632_;
  assign _0466_ = _0364_ | _0109_;
  assign _0661_ = _1687_ | _0103_;
  assign _0020_ = _0649_ | _0648_;
  assign _0712_ = _0151_ | _0116_;
  assign _0851_ = _0386_ | _1688_;
  assign _1689_ = _1690_ | _0361_;
  assign _1691_ = _1692_ | _0197_;
  assign _0298_ = _0177_ | _0269_;
  assign _0762_ = _0529_ | _0267_;
  assign _0736_ = _1694_ | _1693_;
  assign _1079_ = _1695_ | _0615_;
  assign _0773_ = _0250_ | _0552_;
  assign _1402_ = _0195_ | _0607_;
  assign _0764_ = _1696_ | _0748_;
  assign _1286_ = _0228_ | _1033_;
  assign _0940_ = _0338_ | _1697_;
  assign _1698_ = _1203_ | _0270_;
  assign _0345_ = _0144_ | _1374_;
  assign _0272_ = _0232_ | _0290_;
  assign _1549_ = _1699_ | _0171_;
  assign _1429_ = _0042_ | _1700_;
  assign _0792_ = _0213_ | _0144_;
  assign _0883_ = _0042_ | _1024_;
  assign _1132_ = _1701_ | _1567_;
  assign _1233_ = _0097_ | _0255_;
  assign _0728_ = _1304_ | _0345_;
  assign _0559_ = _1206_ | _1028_;
  assign _1702_ = _0489_ | _0102_;
  assign _0553_ = _0615_ | _1703_;
  assign _0004_ = _0209_ | _0406_;
  assign _1704_ = _1686_ | _1028_;
  assign _0778_ = _0857_ | _1705_;
  assign _0779_ = _0619_ | _0635_;
  assign _1513_ = _0456_ | _1211_;
  assign _0461_ = _1707_ | _1706_;
  assign _1708_ = _1709_ | _1348_;
  assign _1711_ = _1712_ | _0879_;
  assign _1138_ = _0065_ | _0625_;
  assign _1453_ = _0930_ | _0134_;
  assign _0437_ = _0356_ | _1713_;
  assign _0898_ = _1088_ | _0488_;
  assign _1436_ = _0069_ | _1645_;
  assign _0075_ = _1527_ | _1019_;
  assign _0812_ = _1714_ | _0193_;
  assign _1528_ = _0208_ | _0059_;
  assign _0219_ = _0304_ | _0463_;
  assign _0871_ = _1715_ | _0452_;
  assign _1206_ = _0019_ | _1716_;
  assign _0362_ = _1464_ | _0357_;
  assign _1203_ = _0058_ | _0993_;
  assign _0487_ = _1064_ | _0271_;
  assign _1199_ = _0071_ | _0914_;
  assign _1238_ = _0088_ | _1718_;
  assign _0881_ = _1691_ | _1719_;
  assign _1720_ = _0134_ | _0893_;
  assign _1172_ = _0214_ | _1056_;
  assign _1721_ = _0566_ | _1046_;
  assign _0383_ = _0226_ | _1551_;
  assign _1722_ = _0091_ | _0263_;
  assign _0855_ = _0708_ | _0909_;
  assign _0141_ = _1716_ | _0197_;
  assign _1723_ = _0195_ | _1724_;
  assign _1725_ = _0241_ | _0613_;
  assign _0539_ = _1048_ | _1102_;
  assign _1654_ = out_data[896] | _0046_;
  assign _1726_ = _0164_ | _0581_;
  assign _1274_ = _1728_ | _1727_;
  assign _1729_ = _0019_ | _1730_;
  assign _0999_ = _0096_ | _0103_;
  assign _0127_ = _0189_ | _0250_;
  assign _0882_ = _1654_ | _0613_;
  assign _1580_ = _0325_ | _0032_;
  assign _0069_ = _0524_ | _0609_;
  assign _1166_ = _1247_ | _0780_;
  assign _0569_ = _0677_ | _1733_;
  assign _1734_ = _0454_ | _0299_;
  assign _1221_ = _0835_ | _0620_;
  assign _1294_ = _1735_ | _0206_;
  assign _1737_ = _0134_ | _1421_;
  assign _1136_ = _0999_ | _0134_;
  assign _0118_ = in_data[1671] | _0401_;
  assign _1204_ = _1738_ | _0226_;
  assign _1739_ = _1740_ | _0466_;
  assign _1258_ = _0151_ | _0337_;
  assign _1741_ = _0873_ | _0730_;
  assign _1742_ = _0145_ | _0420_;
  assign _1176_ = _0027_ | _1072_;
  assign _1744_ = _1004_ | _0367_;
  assign _1192_ = _1745_ | _0192_;
  assign _0980_ = _0721_ | _0426_;
  assign _0136_ = _0128_ | _1747_;
  assign _1606_ = _0053_ | _0663_;
  assign _1603_ = _0753_ | _0082_;
  assign _1198_ = _0462_ | _1749_;
  assign _1752_ = _0669_ | _0623_;
  assign _1310_ = _0343_ | _0025_;
  assign _0021_ = _1753_ | _0042_;
  assign _0531_ = _0025_ | _0311_;
  assign _1758_ = _1759_ | _1691_;
  assign _1760_ = _0171_ | _1761_;
  assign _0152_ = _0189_ | _1755_;
  assign _0174_ = _0320_ | _0265_;
  assign _0924_ = _0739_ | _0603_;
  assign _0453_ = _1768_ ^ _1690_;
  assign _0099_ = _1000_ ^ _0116_;
  assign _0017_ = _1134_ ^ _0800_;
  assign _0748_ = _1771_ ^ _0134_;
  assign _1772_ = _1540_ ^ _0416_;
  assign _0087_ = _0191_ ^ _0517_;
  assign _1777_ = _0439_ ^ _0590_;
  assign _1655_ = _0678_ ^ _0118_;
  assign _0615_ = _0162_ ^ _0490_;
  assign _1780_ = _0336_ ^ _0055_;
  assign _0983_ = _0193_ ^ _0134_;
  assign _0368_ = _0238_ ^ _0609_;
  assign out_data[1504] = _0959_ ^ _1621_;
  assign out_data[1376] = _1783_ ^ _1782_;
  assign out_data[928] = _0707_ ^ _0566_;
  assign out_data[512] = _1784_ ^ _0196_;
  assign out_data[448] = _1370_ ^ _0955_;
  assign out_data[0] = _0117_ ^ _0465_;
  assign _0194_ = _0189_ ^ _0154_;
  assign _0132_ = _0277_ ^ _0103_;
  assign _1000_ = _1785_ ^ _0025_;
  assign _0160_ = _0334_ ^ _1786_;
  assign _0697_ = _0857_ ^ _0769_;
  assign _0891_ = _0099_ ^ _0566_;
  assign _1750_ = _0318_ ^ _0315_;
  assign _0175_ = _0587_ ^ _0633_;
  assign _0690_ = _1787_ ^ _0226_;
  assign _0024_ = _0856_ ^ _0152_;
  assign _0645_ = _1788_ ^ _0043_;
  assign _0258_ = _0096_ ^ _0043_;
  assign _0994_ = _1790_ ^ _1789_;
  assign _0420_ = _1791_ ^ out_data[416];
  assign _0620_ = _1792_ ^ _0924_;
  assign _0149_ = _1793_ ^ _0082_;
  assign _0023_ = _0043_ ^ _0024_;
  assign _0235_ = _0438_ ^ _0134_;
  assign _1483_ = _0129_ ^ _1794_;
  assign _0281_ = _0318_ ^ _0294_;
  assign _0009_ = _1795_ ^ _0016_;
  assign _1368_ = _0067_ ^ _0506_;
  assign _1348_ = _1064_ ^ _0228_;
  assign _0452_ = _0661_ ^ _0185_;
  assign _0450_ = _0105_ ^ _0128_;
  assign _0317_ = _0103_ ^ _1000_;
  assign _1265_ = _0315_ ^ _0857_;
  assign _1464_ = _0566_ ^ _0151_;
  assign _1552_ = _0071_ ^ _0454_;
  assign _0656_ = _1797_ ^ _1796_;
  assign _1072_ = _0270_ ^ _0204_;
  assign _1561_ = _0203_ ^ _0325_;
  assign _1211_ = _0127_ ^ _0404_;
  assign _1550_ = _1798_ ^ _1134_;
  assign _0012_ = _0197_ ^ _0620_;
  assign _1343_ = _0581_ ^ _0303_;
  assign _0899_ = _0617_ ^ _0290_;
  assign _1634_ = _0608_ ^ _1086_;
  assign _1799_ = _1348_ ^ _1551_;
  assign _0755_ = _0611_ ^ _0035_;
  assign _0275_ = _1800_ ^ _0359_;
  assign _0649_ = _0228_ ^ _0309_;
  assign _0585_ = _1801_ ^ _0128_;
  assign _0979_ = _0092_ ^ _0343_;
  assign _0722_ = _0014_ ^ _0158_;
  assign _0939_ = _0419_ ^ _1170_;
  assign _0287_ = _1804_ ^ _1803_;
  assign _0264_ = _1805_ ^ _0134_;
  assign _1379_ = _1806_ ^ _0170_;
  assign _0949_ = _1807_ ^ _0593_;
  assign _1645_ = _0615_ ^ _0700_;
  assign _0550_ = _0999_ ^ _0193_;
  assign _0337_ = _1024_ ^ _0626_;
  assign _1059_ = _1621_ ^ _1750_;
  assign _1147_ = _0071_ ^ _0200_;
  assign _1808_ = _0259_ ^ _0730_;
  assign _1447_ = _0211_ ^ _0463_;
  assign _1809_ = _0401_ ^ _1265_;
  assign _0458_ = _0194_ ^ _0019_;
  assign _0106_ = _0993_ ^ _0125_;
  assign _0314_ = _0140_ ^ _0317_;
  assign _0519_ = _0258_ ^ _1810_;
  assign _0711_ = _0752_ ^ _0071_;
  assign _1195_ = _1352_ ^ _1811_;
  assign _1812_ = _0166_ ^ _1128_;
  assign _0561_ = _1813_ ^ _0535_;
  assign _0031_ = _1814_ ^ _0519_;
  assign _0048_ = _0997_ ^ _0706_;
  assign _1093_ = _0097_ ^ _1034_;
  assign _0787_ = _1815_ ^ _0194_;
  assign _0580_ = _1816_ ^ _0259_;
  assign _1099_ = _1817_ ^ _0041_;
  assign _0523_ = _0651_ ^ _1393_;
  assign _0849_ = _1096_ ^ _0042_;
  assign _0578_ = _0376_ ^ _0687_;
  assign _0946_ = _0148_ ^ _1461_;
  assign _0241_ = in_data[2079] ^ in_data[554];
  assign _1818_ = _0573_ ^ _0532_;
  assign _0944_ = _0595_ ^ _1598_;
  assign _1405_ = _0056_ ^ _0620_;
  assign _1421_ = _0458_ ^ _1047_;
  assign _0708_ = _0565_ ^ _0103_;
  assign _1182_ = _0680_ ^ _0159_;
  assign _0121_ = _0228_ ^ _0205_;
  assign _1820_ = _1683_ ^ _0811_;
  assign _1179_ = _0354_ ^ _0117_;
  assign _1602_ = _1821_ ^ _1474_;
  assign _0151_ = _0320_ ^ _0638_;
  assign _1231_ = _1348_ ^ _0140_;
  assign _1822_ = _0609_ ^ _0591_;
  assign _1090_ = _1705_ ^ _0828_;
  assign _0373_ = _0116_ ^ _1669_;
  assign _1733_ = _0144_ ^ _0612_;
  assign _1251_ = _0481_ ^ _0891_;
  assign _1472_ = _0314_ ^ _0193_;
  assign _0900_ = _0469_ ^ _0117_;
  assign _0930_ = _1820_ ^ _1824_;
  assign _1298_ = _0151_ ^ _1825_;
  assign _0325_ = _1506_ ^ _0071_;
  assign _1718_ = _0338_ ^ _0949_;
  assign _1551_ = _0189_ ^ _0524_;
  assign _1746_ = _0232_ ^ _1018_;
  assign _1827_ = _0175_ ^ _1738_;
  assign _1456_ = _0108_ ^ _0259_;
  assign _1505_ = _0848_ ^ _0141_;
  assign _1828_ = _0697_ ^ _1829_;
  assign _0061_ = _1702_ ^ _0598_;
  assign _0956_ = _1830_ ^ _0481_;
  assign _1831_ = _1303_ ^ _1134_;
  assign _1832_ = _0348_ ^ _0453_;
  assign _0576_ = _0656_ ^ _1833_;
  assign _1834_ = _0221_ ^ _0891_;
  assign _0958_ = _1336_ ^ _0219_;
  assign _0334_ = _1551_ ^ _0317_;
  assign _0825_ = _0234_ ^ _0214_;
  assign _1835_ = _1655_ ^ _0348_;
  assign _0028_ = _0700_ ^ _0149_;
  assign _0177_ = _0287_ ^ _0082_;
  assign _0462_ = _0015_ ^ _1836_;
  assign _0948_ = _1837_ ^ _0061_;
  assign _1117_ = _0851_ ^ _1838_;
  assign _0457_ = _0712_ ^ _1839_;
  assign _1124_ = _0096_ ^ _1112_;
  assign _0625_ = _0270_ ^ _0401_;
  assign _1841_ = _0102_ ^ _0727_;
  assign _0971_ = _0565_ ^ _1031_;
  assign _1614_ = _0225_ ^ _0099_;
  assign _0817_ = _0747_ ^ _0134_;
  assign _1500_ = _1061_ ^ _1318_;
  assign _0424_ = _0774_ ^ _0032_;
  assign _1843_ = _0454_ ^ _0146_;
  assign _0440_ = _0708_ ^ _1844_;
  assign _1845_ = _0025_ ^ _0209_;
  assign _0942_ = _1266_ ^ _0058_;
  assign _1292_ = _1290_ ^ _1027_;
  assign _0431_ = _1846_ ^ _0039_;
  assign _1847_ = _0401_ ^ _1848_;
  assign _0872_ = _1703_ ^ _1850_;
  assign _1852_ = _0341_ ^ _0068_;
  assign _0868_ = _0227_ ^ _1518_;
  assign _0511_ = _1046_ ^ _0355_;
  assign _1540_ = _0812_ ^ _0298_;
  assign _1595_ = _1854_ ^ _0732_;
  assign _1533_ = _0413_ ^ _1595_;
  assign _0893_ = _0151_ ^ _1307_;
  assign _1858_ = _0384_ ^ _1859_;
  assign _0054_ = _1861_ ^ _0697_;
  assign _1862_ = _1258_ ^ _0261_;
  assign _1863_ = _0664_ ^ _1718_;
  assign _0111_ = _0043_ ^ _1511_;
  assign _1864_ = _1741_ ^ _0462_;
  assign _0589_ = _0146_ ^ _0071_;
  assign _1865_ = _0682_ ^ _1056_;
  assign _0065_ = _0144_ ^ _0318_;
  assign _1867_ = _1089_ ^ _1799_;
  assign _1868_ = _0065_ ^ _1129_;
  assign _0544_ = _1869_ ^ _1867_;
  assign _1626_ = _0103_ ^ _0475_;
  assign _0074_ = _1549_ ^ _0046_;
  assign _1607_ = _0234_ ^ _0014_;
  assign _1870_ = _0748_ ^ _0831_;
  assign _1209_ = _0489_ ^ _1454_;
  assign _1784_ = _0643_ ^ _1514_;
  assign _1873_ = _1084_ ^ _0639_;
  assign _0546_ = _0449_ ^ _1874_;
  assign _0912_ = _0562_ ^ _1875_;
  assign _0014_ = _0101_ ^ _0022_;
  assign _1876_ = _1483_ ^ _0900_;
  assign _1878_ = _1879_ ^ _0875_;
  assign _1880_ = _1208_ ^ _0094_;
  assign out_data[64] = _1881_ ^ _0957_;
  assign _1009_ = _0227_ ^ _0226_;
  assign _1883_ = _0032_ ^ _0144_;
  assign _1884_ = _0196_ ^ _1885_;
  assign { _0596_, _1753_, _1889_[10:8], _1624_, _1312_, _1889_[5:0] } = { _1891_[12:5], _0639_, _1009_, _0109_, _1283_, _0219_ } + { _0588_, _1890_[11], _0350_, _0716_, _1890_[8:6], _1136_, _0238_, _0109_, _0306_, _0116_, _0238_ };
  assign _1892_ = { _1894_[55:48], _0043_, _0213_, _1894_[45:41], _0676_, _1894_[39:38], _0445_, _0179_, _0496_, _0476_, _0054_, _0677_, _0349_, _1025_, _0298_, _1171_, _1218_, _0269_, _0476_, _0470_, _1733_, _1065_, _0390_, _1220_, _0886_, _1894_[18:3], _0043_, _0944_, _0076_ } + { _0766_, _0490_, _0526_, _1609_, _0241_, _1893_[50:49], _0771_, _0807_, _0894_, _0551_, _1893_[44:14], _0702_, _1402_, _1153_, _1893_[10:7], _1034_, _1893_[5:4], _1374_, _1787_, _0126_, _1328_ };
  assign { _1897_[53:52], _1665_, _1897_[50:27], _1260_, _1897_[25:21], _0037_, _1897_[19:0] } = { _1899_[53:3], _0079_, _0911_, _0303_ } + { _0405_, _0922_, _0062_, _1036_, _0381_, _0289_, _0636_, _0565_, _0398_, _1182_, _0884_, _0526_, _0599_, _1171_, _0858_, _1898_[38:23], _1517_, _1898_[21:17], _1593_, _1898_[15:10], _0765_, _1898_[8:0] };
  assign { _1902_[38:29], _1293_, _1902_[27:0] } = { _1904_[38:22], _1599_, _1893_[44:38], _0698_, _0821_, _1812_, _0971_, _1904_[9:2], _0272_, _0001_ } + { _1903_[38:36], _1213_, _1903_[34:3], _1742_, _1555_, _1149_ };
  assign { _0077_, _1905_[3:0] } = { _1906_[4:1], _0744_ } + { _1890_[11], _0350_, _0935_, _0493_, _1852_ };
  assign { _1918_[31:11], _1295_, _1918_[9:2], _0937_, _1918_[0] } = { _1920_[31:22], _0056_, _1920_[20:19], _1816_, _1920_[17:16], _1168_, _1920_[14:2], _1841_, _0299_ } + { _1919_[31:17], _0557_, _1919_[15:7], _1882_, _1919_[5], _0904_, _1125_, _1025_, _0882_, _0856_ };
  assign out_data[1997:1984] = { _0764_, _0206_, _1947_[11:6], _1267_, _1947_[4:3], _1646_, _0522_, _0149_ } + { _1946_[13:1], _1462_ };
  assign out_data[1417:1408] = { _1949_[9:5], _1883_, _0366_, _0372_, _0982_, _0025_ } + _1948_;
  assign { _1950_[215:196], out_data[1311:1280], _1950_[163:0] } = { _1952_[215:214], _1083_, _1952_[212:206], _1246_, _1952_[204:184], _1389_, _1952_[182:177], _0344_, _1952_[175:165], _1194_, _1952_[163:157], _0228_, _1758_, _1659_, _0292_, _0054_, _1144_, _1777_, _0420_, _0357_, _0145_, _0044_, _0701_, _1021_, _0804_, _1014_, _1952_[141], _1621_, _1577_, _1320_, _1952_[137], _1648_, _0278_, _0811_, _0855_, _1657_, _0028_, _1780_, _0683_, _1362_, _0175_, _1301_, _0029_, _1433_, _1177_, _1138_, _0797_, _1892_, _0939_, _0362_, _0324_, _0379_, _1215_, _1952_[59:45], _1232_, _1494_, _1952_[42], _0803_, _1952_[40:17], _1586_, _1952_[15:12], _1385_, _1952_[10:7], _1118_, _1952_[5:4], out_data[1888], _1554_, _0217_, _1044_ } + { _1897_[47:27], _1260_, _1897_[25:21], _0037_, _1897_[19:4], _0228_, _0625_, _1951_[169:159], _1255_, _1951_[157:151], _1276_, _1951_[149:144], _1042_, _1951_[142:139], _0124_, _0929_, _1951_[136:134], _0505_, _0423_, _0087_, _1951_[130:128], _0235_, _0917_, _0917_, out_data[544], _1951_[123], _1122_, _1951_[121:119], _1609_, _0080_, _1951_[116:105], _1560_, _1951_[103:88], _1910_[9:3], _1951_[80:58], _0285_, _0868_, _0977_, _1429_, _0413_, _0879_, _1486_, _0334_, _0032_, _0412_, _0118_, _1085_, _0529_, _0217_, _1880_, _0442_, _0325_, _1178_, _0015_, _1561_, _0964_, _1831_, _1555_, _1606_, _1951_[33], _1412_, _1951_[31], _1496_, _1951_[29:6], _0382_, _1951_[4:2], _0800_, _1371_ };
  assign out_data[1276:1248] = { _1954_[28:12], _1872_, _1954_[10:9], out_data[1952], _1954_[7:0] } + { _1935_[75:72], _1953_[24:8], _1428_, _1953_[6], _0611_, _1463_, _0835_, _1033_, _1599_, _1664_ };
  assign out_data[1150:1120] = { _1956_[30:24], _1618_, _1956_[22], _1642_, _1629_, _0017_, _1956_[18:15], _0506_, _1956_[13:12], _0828_, _1956_[10:2], _0218_, _0273_ } + { _1952_[52:48], _1955_[25:20], _0072_, _1955_[18], _1853_, _1955_[16], _1487_, _1955_[14:1], _0217_ };
  assign out_data[1101:1088] = { _1958_[13:4], _0661_, _0875_, _0359_, _1137_ } + { _1904_[36:31], _0950_, _1190_, _0933_, _0358_, _0102_, _1870_, _1957_[1:0] };
  assign out_data[809:800] = { _0633_, _0162_, _1959_[7], _1202_, _1431_, _1959_[4:3], _1145_, _1089_, _0948_ } + { _0760_, _1901_[12:10], _0879_, _1901_[8:6], _0533_, out_data[960] };
  assign { out_data[639:608], _1960_[2:0] } = { out_data[1276:1254], _1962_[11:5], _1261_, _1962_[3:1], _0228_ } + { _1961_[34:1], _0000_ };
  assign { _1963_[76:60], out_data[511:480], _1963_[27:0] } = { _1950_[152:87], _0071_, _0727_, _1289_, _0881_, _0816_, _0166_, out_data[1664], _1574_, _0876_, _0194_, _0760_ } + { _1452_, _1964_[75:74], _1647_, _1964_[72:67], _0364_, _1888_[13], _0036_, _0706_, _1888_[10:5], _0673_, _1964_[55], _1679_, _1617_, _1964_[52], _1795_, _1964_[50:48], _1016_, _1964_[46:45], _0492_, _1964_[43], _1706_, _0890_, _1084_, _1831_, _0843_, _0721_, _0960_, _0480_, _0268_, _1381_, _1964_[32:31], _1156_, _1964_[29:27], _1264_, _1299_, _0568_, _0915_, _0355_, _1964_[21:7], _1092_, _0232_, _0615_, out_data[864], _0934_, _0018_, _1394_ };
  assign { out_data[319:288], _1965_[45:0] } = { _1920_[16], _1168_, _1920_[14], _0241_, _0752_, _1079_, _0756_, _0082_, _0586_, _1063_, _0025_, _1913_[36:31], _1466_, _1913_[29:25], _0567_, _1701_, _1913_[22:10], _1821_, _1913_[8], _1259_, _0301_, _1967_[35:23], _1123_, _1967_[21:15], _1668_, _1967_[13:10], _1321_, _0473_, _1967_[7:0] } + { _1966_[77:65], _1052_, _0447_, _0096_, _1275_, _1299_, _0062_, _1207_, _1580_, _1876_, _0189_, _0068_, _1043_, _1933_[13:9], _1244_, _1933_[7:6], _1966_[44:42], _1236_, _1174_, _1966_[39:34], _0990_, _1966_[32:27], _0988_, _1879_, _1966_[24:19], _0528_, _1966_[17:14], _0540_, _1864_, _1186_, _1505_, _1966_[9], _0631_, _1744_, _0259_, _1549_, _1966_[4], _0818_, _1966_[2], _0807_, _0636_ };
  assign { _0719_, _1968_[50], _1022_, _1968_[48:14], _0142_, _1968_[12:0] } = { _1970_[51:20], _1253_, _1970_[18:16], _1210_, _1682_, _1970_[13:11], _0159_, _1786_, _0402_, _1397_, _1569_, _1970_[5], _0716_, _0907_, _0206_, _0241_, _0071_ } + { _1969_[51:36], _0677_, _1969_[34:29], _0985_, _1969_[27:8], _0453_, _1266_, _0096_, _0529_, _0752_, _1283_, _0625_, _0065_ };
  assign { _1971_[25:19], _0922_, _1971_[17:13], _1525_, _1971_[11:0] } = { _1973_[25:24], _0504_, _1597_, _0684_, _1973_[20:19], _1970_[51:39], _0464_, _1235_, _1374_, _0356_, _0999_, _0194_ } + { _1972_[25:22], _1687_, _1972_[20:11], _1310_, _0636_, _0678_, _0993_, _0403_, _0589_, _0739_, _0918_, _0101_, _0639_, _0518_ };
  assign { _0155_, _1974_[0] } = { _0356_, _0733_ } + { _0059_, _0205_ };
  assign { _1975_[74:54], _1790_, _1975_[52], _1926_[30:5], _0614_, _1926_[3:2], _1975_[22:0] } = { _1889_[2], _1976_[70:58], _1797_, _1976_[56:34], _0100_, _1976_[32:26], _1341_, _1976_[24:23], _1977_[25:24], _1243_, _1384_, _1669_, _0256_, _0116_, _1203_, _0983_, _1046_, _0915_, _0019_, _0227_, _0356_, _1621_, _0155_, _1974_[0], _1527_, _1374_, _0217_, _0043_, _0134_, _0069_, _0311_, _0134_, _0046_ } + { _0189_, _0033_, _0065_, _0018_, _1976_[70:58], _1797_, _1976_[56:34], _0100_, _1976_[32:26], _1341_, _1976_[24:23], _0121_, _0563_, _0591_, _1976_[19:16], _1335_, _1976_[14], _0172_, _0120_, _1568_, _1976_[10:9], _0604_, _1976_[7], _0945_, _1976_[5], _0602_, _1976_[3:0] };
  assign { _1978_[58:49], _1446_, _1940_[36:26], _1696_, _1940_[24], _1230_, _1940_[22:20], _1901_[86:74], _0107_, _1901_[72:70], _1978_[13:0] } = { _1976_[37:36], _1979_[56:55], _1658_, _1979_[53], _1268_, _1979_[51:43], _1002_, _1979_[41:22], _0790_, _1979_[20:16], _1562_, _1979_[14:9], _1616_, _1979_[7], _1621_, _0238_, _0071_, _0401_, _0287_, _0857_, _0049_ } + { _1968_[45:14], _0142_, _1968_[12:9], _1964_[67], _0364_, _1888_[13], _0036_, _0706_, _1888_[10:5], _0673_, _1964_[55], _1679_, _0361_, _0401_, _0174_, _0200_, _0159_, _0287_, _0272_, _0609_ };
  assign { _1956_[18:15], _0506_, _1956_[13:12] } = { _0293_, _0082_, _0490_, _0563_, _0118_, _0250_, _0154_ } + { in_data[1353:1349], _0317_, _0320_ };
  assign { _0993_, _0403_ } = { _0200_, _0573_ } + { _0529_, _0103_ };
  assign { _1980_[23:6], _1367_, _1980_[4], _1681_, _1980_[2:0] } = { _1381_, _1520_, _1982_[21:16], _1534_, _1982_[14:6], _1287_, _0174_, _0343_, _0383_, _0265_, _0453_ } + { _0025_, _0238_, _0617_, _0625_, _0025_, _0151_, _0043_, _0469_, _1951_[33], _1412_, _1951_[31], _1496_, _1981_[11:9], _0299_, _0223_, _1981_[6:2], _1794_, _0194_ };
  assign { _1983_[46:26], _1928_[24:18], _0244_, _1928_[16:12], _0441_, _1928_[10:9], _1983_[9:0] } = { _1984_[46:39], _1714_, _1984_[37:36], _0251_, _1984_[34:15], _0243_, _0739_, _1153_, _1893_[10:7], _1034_, _1893_[5:4], _1374_, _1787_, _0126_, _1328_, _0254_ } + { _1969_[45:36], _0677_, _1969_[34:29], _0985_, _1969_[27:14], _0594_, _0097_, _0615_, _0587_, _0174_, _1205_, _1810_, _0123_, _1932_[6], _0595_, _0096_, _0238_, _0098_, _0250_, _0154_ };
  assign { _1985_[11:2], _1692_, _1985_[0] } = { _0350_, _0716_, _0565_, _0572_, _1374_, _1527_, _0518_, _1225_, _1141_, _0622_, _1986_[1], _0068_ } + { _1786_, _0402_, _1397_, _1569_, _1970_[5], _0206_, _0316_, _0097_, _0936_, _0566_, _0287_, _0265_ };
  assign { _1987_[54:52], _1596_, _1987_[50:48], _1839_, _1987_[46:31], _0693_, _1987_[29:23], _0798_, _1987_[21:0] } = { _1989_[54:33], _1344_, _1989_[31:5], _1792_, _1989_[3:2], _0134_, _0311_ } + { _1988_[54:51], _0291_, _1988_[49], _1383_, _1988_[47:46], _1697_, _1988_[44:43], _0277_, _1988_[41:38], _0130_, _1988_[36], _0725_, _1988_[34:27], _1406_, _1175_, _1988_[24], _0921_, _1988_[22], _1819_, _1988_[20:19], _0102_, _0697_, _0690_, _1964_[67], _0364_, _1888_[13], _0036_, _0706_, _1888_[10:5], _0673_, _1964_[55], _1679_, _0589_, _0096_ };
  assign { _1990_[55], _1811_, _1990_[53], _1413_, _1990_[51:45], _1764_, _1990_[43:23], _1074_, _1990_[21:16], _0928_, _1990_[14:13], _0495_, _1990_[11:0] } = { _1989_[48:33], _1344_, _1989_[31:5], _1792_, _1989_[3:2], _1992_[8], _0189_, _0221_, _0566_, _1992_[4:0] } + { _1991_[55:47], _1193_, _1553_, _1991_[44:43], _0219_, _0887_, _0359_, _0642_, _0019_, _1951_[169:159], _1255_, _1951_[157:151], _1276_, _1951_[149:144], _1042_, _1951_[142:139], _0124_, _0929_, _1951_[136:134], _0678_, _1007_ };
  assign { _1993_[9:6], _1041_, _1993_[4:0] } = { _1994_[9:6], _0840_, _1994_[4:3], _0597_, _0594_, _0999_ } + { _1900_[70], _0389_, _1900_[68:66], _0833_, _1305_, _1900_[63], _0096_, _0325_ };
  assign { _1995_[17:14], _0224_, _1995_[12:6], _1242_, _1995_[4:1], _1011_ } = { _1969_[22:9], _0136_, _0565_, _0043_, _0057_ } + { in_data[836:826], _1203_, _1716_, _1996_[4], _1365_, _0104_, _1476_, _1467_ };
  assign { _1966_[4], _0818_, _1966_[2] } = { _0581_, _0092_, _0160_ } + _1997_;
  assign { _1998_[40:30], _1325_, _1998_[28:0] } = { _1976_[64:58], _1797_, _1976_[56:34], _0100_, _1976_[32:26], _1341_, _1976_[24] } + in_data[1270:1230];
  assign { _1999_[139:120], _1109_, _1999_[118:100], _1030_, _1999_[98:76], _1817_, _1999_[74:67], _0574_, _1999_[65:32], _1303_, _1999_[30:0] } = { _2001_[139:138], _0211_, _2001_[136:113], _0752_, _2001_[111], _1323_, _2001_[109], _1309_, _1081_, _2001_[106:103], _1351_, _2001_[101:99], _1353_, _2001_[97], _1359_, _2001_[95:86], _0998_, _2001_[84:73], _1765_, _2001_[71], _0719_, _1968_[50], _1022_, _1968_[48:14], _0142_, _1968_[12:0], _0287_, _0290_, _0015_, _0368_, _0278_, _0434_, _1985_[11:2], _1692_, _1985_[0], _0521_ } + { _1908_[10], _0535_, _1908_[8:7], _0363_, _0325_, _0210_, _0155_, _1974_[0], _0566_, _1007_, _0096_, _1951_[33], _1412_, _1951_[31], _1496_, _2000_[123:108], _1361_, _2000_[106:100], _1506_, _2000_[98], _0113_, _2000_[96:92], _0313_, _2000_[90:86], _0737_, _2000_[84:80], _0401_, _0105_, _0082_, _0152_, _0642_, _0108_, _0572_, _0317_, _0057_, _1951_[33], _1412_, _1951_[31], _1496_, _1225_, _1141_, _0622_, _1986_[1], _0095_, _1393_, _0241_, _2000_[59:50], _1570_, _2000_[48:46], _1314_, _1419_, _0391_, _2000_[42:35], _1747_, _2000_[33:31], _1307_, _2000_[29:27], _1318_, _0097_, _1009_, _0502_, _0401_, _0125_, _2000_[20:19], _0564_, _2000_[17:14], _0925_, _1939_[12:8], _0501_, _1939_[6], _1306_, _2000_[4:3], _1632_, _1373_, _2000_[0] };
  assign { _2003_[10:9], _1126_, _1631_, _2003_[6:3], _1372_, _1217_, _2003_[0] } = { _2005_[10:8], _1327_, _2005_[6:4], _0189_, _0320_, _0278_, _0988_ } + { _2004_[10:6], _1387_, _0581_, _0572_, _0318_, _0359_, _0117_ };
  assign { _1677_, _0409_, _1804_, _1386_, _2002_[27:26], _1381_, _1520_, _1982_[21:16], _1534_, _1982_[14:6], _1287_, _2002_[6:0] } = { _0132_, _0068_, _0043_, _0356_, _0238_, _0189_, _0103_, _1153_, _1893_[10:7], _1034_, _1893_[5:4], _1374_, _1787_, _0126_, _1328_, _0241_, _1153_, _1893_[10:7], _1034_, _1893_[5:4], _1374_, _1787_, _0126_, _1328_ } + { in_data[1485:1473], _1153_, _1893_[10:7], _1034_, _1893_[5:4], _1374_, _1787_, _0126_, _1328_, _0128_, _0277_, _0127_, _0128_, _0082_, _0238_, _0189_ };
  assign { _1254_, _0468_, _2006_[6], _0404_, _2006_[4:3], _1931_[3], _1308_, _0513_ } = { _0993_, _0359_, _0134_, _0103_, _0132_, _0025_, _0356_, _0277_, _0359_ } + { _2007_[8:1], _0103_ };
  assign { _2008_[14:3], _1531_, _1068_, _2008_[0] } = { _1952_[209:206], _1246_, _1952_[204:196], _0221_ } + { _1386_, _2002_[27:26], _1381_, _1520_, _1982_[21:16], _1534_, _1982_[14:13], _0277_ };
  assign { _1805_, _2009_[2], _0819_, _1807_ } = { _0343_, _0135_, _1205_, _0152_ } + { _2010_[3:1], _0240_ };
  assign { _2011_[43:28], _1044_, _2011_[26:6], _0181_, _2011_[4:0] } = { _2012_[43:28], _1625_, _2012_[26:22], _1678_, _1222_, _2012_[19:2], _1613_, _0082_ } + { _1596_, _1987_[50:48], _1839_, _1987_[46:31], _0693_, _1987_[29:23], _0798_, _1987_[21:8] };
  assign { _2013_[17:10], _1857_, _2013_[8:7], _1829_, _1040_, _2013_[4:0] } = { _2014_[17:10], _1988_[54:51], _0291_, _1988_[49], _1383_, _1988_[47:46], _0097_ } + { _1990_[27], _2008_[14:3], _1531_, _1068_, _2008_[0], _0529_, _0043_ };
  assign { _0548_, _2015_[20:2], _1369_, _2015_[0] } = { _2000_[20:19], _0564_, _2000_[17:14], _0925_, _1939_[12:8], _0501_, _1939_[6], _1306_, _2000_[4:3], _1632_, _1373_, _0609_, _0137_ } + { _2016_[21:6], _0145_, _0122_, _0042_, _1449_, _0594_, _0781_ };
  assign { _2017_[65:61], _1364_, _2017_[59:37], _1410_, _2017_[35:33], _0414_, _2017_[31:14], _1442_, _2017_[12:0] } = { _1970_[42:38], _0117_, _0272_, _2019_[58:57], _1636_, _2019_[55:37], _0070_, _1920_[31:22], _0056_, _1920_[20:19], _1816_, _1920_[17:16], _1168_, _1920_[14:2], _2019_[5], _1655_, _0452_, _0095_, _0318_, _0873_ } + { _0920_, _2004_[10:6], _1387_, _2018_[58:56], _0397_, _1640_, _2018_[53], _0023_, _1449_, _0191_, _1265_, _0589_, _0907_, _0620_, _0206_, _0311_, _2000_[20:19], _0564_, _2000_[17:14], _0925_, _1939_[12:8], _0501_, _1939_[6], _1306_, _2000_[4:3], _1632_, _1373_, _2000_[0], _0795_, _0108_, _1203_, _0854_, _0986_, _1908_[14:13], _1564_, _1908_[11:10], _0535_, _1908_[8:7], _0984_, _0477_, _1329_, _0716_, _0600_, _0146_, _0572_, _0856_, _0134_, _0692_ };
  assign { _1912_[29:15], _1592_, _1912_[13:10], _0188_, _1912_[8:2] } = { in_data[1421:1397], _0311_, _0678_, _0348_ } + { _1985_[5:2], _1692_, _0235_, _0275_, _0316_, _0272_, _0325_, _1046_, _0324_, _1322_, _0254_, _0469_, _0044_, _1493_, _2020_[10:9], _0293_, _2020_[7:5], _0044_, _0608_, _0178_, _0726_, _0715_ };
  assign { _1909_[12], _1908_[39:38], _1885_, _1908_[36], _1270_, _1908_[34], _1048_, _1909_[4:2], _1167_ } = _1943_[102:91] + { _2013_[8:7], _1829_, _1040_, _2013_[4:2], _0270_, _0043_, _0122_, _0068_, _0581_ };
  assign { _2021_[21:18], _0688_, _2021_[16:13], _1189_, _2021_[11:0] } = { _0208_, _0235_, _0986_, _1908_[14:13], _1564_, _1908_[11:10], _0535_, _1908_[8:7], _1561_, _0619_, _2022_[8:6], _1160_, _2022_[4:3], _1069_, _2022_[1:0] } + { _1952_[189:184], _1389_, _1952_[182:177], _0344_, _1952_[175:169], _0626_ };
  assign { _2023_[13:12], _1469_, _1408_, _2023_[9:7], _0327_, _2023_[5:0] } = { _2024_[13:12], _1825_, _2024_[10:2], _0274_, _0016_ } + { _1990_[13], _0495_, _1909_[12], _1908_[39:38], _1885_, _1908_[36], _1270_, _1908_[34], _1048_, _1909_[4:2], _1167_ };
  assign { _1952_[59:45], _1232_, _1494_, _1952_[42], _0803_, _1952_[40:17], _1586_ } = { _2026_[43:34], _0842_, _2026_[32:11], _1097_, _2026_[9:7], _0116_, _0097_, _1621_, _0111_, _0221_, _0176_, _0309_ } + { _2025_[43:40], _1785_, _2025_[38:34], _1510_, _2025_[32:27], _0896_, _2025_[25], _0290_, _0133_, _0627_, _0043_, _0656_, _0716_, _0145_, _0752_, _1993_[9:6], _1041_, _1993_[4:0], _0627_, _0057_, _0383_, _0620_, _0281_, _0259_, _0058_ };
  assign { _2027_[10:9], _0889_, _2027_[7:5], _0260_, _2027_[3:1], _1107_ } = { _2000_[123:122], _0690_, _1283_, _1077_, _0248_, _1684_, _2028_[3], _1326_, _2028_[1], _0489_ } + _1998_[10:0];
  assign { _1801_, _2029_[42:30], _1012_, _2029_[28:19], _1357_, _2029_[17], _1440_, _2029_[15:11], _1115_, _2029_[9:0] } = { _1999_[57:32], _1303_, _1999_[30:18], _0620_, _0134_, _0317_, _0217_ } + { _1952_[56:45], _1232_, _1494_, _1952_[42], _0803_, _1952_[40:25], _1966_[4], _0818_, _1966_[2], _0357_, _0988_, _1322_, _0152_, _1655_, _1009_, _0258_, _0043_, _0178_ };
  assign { _2030_[66:46], _0705_, _2030_[44:42], _1598_, _2030_[40:16], _1685_, _2030_[14:0] } = { _2032_[66:54], _1527_, _0228_, _0149_, _1265_, _0272_, _0915_, _2008_[14:3], _1531_, _1068_, _2008_[0], _1028_, _2032_[31:26], _1826_, _2032_[24:13], _0606_, _2032_[11:10], _1754_, _2032_[8:1], _0617_ } + { _2031_[66], _0328_, _2031_[64], _0007_, _1699_, _2031_[61:55], _1806_, _2031_[53], _0206_, _2031_[51], _1800_, _2031_[49:47], _1991_[55:47], _1193_, _1553_, _1991_[44:43], _2031_[33:31], _1788_, _2031_[29:23], _0514_, _2031_[21:19], _1887_[16], _2031_[17], _1101_, _1814_, _2031_[14:3], _1509_, _0401_, _0235_ };
  assign { _2033_[23:22], _1783_, _2033_[20:6], _1407_, _2033_[4:0] } = { _2035_[23:19], _1455_, _1507_, _2035_[16], _1674_, _2035_[14:2], _0320_, _0795_ } + { _2034_[23:15], _0000_, _0700_, _0153_, _0634_, _0739_, _0185_, _0146_, _0304_, _0278_, _0238_, _0697_, _0196_, _0589_, _0572_, _0529_ };
  assign { _2036_[16:14], _0509_, _0236_, _2036_[11:3], _1715_, _2036_[1:0] } = { _1995_[15:14], _0224_, _1995_[12:6], _1242_, _1995_[4:1], _1011_, _0175_ } + { _2022_[6], _1160_, _0841_, _0071_, _0166_, _0227_, _1981_[11:9], _0299_, _0223_, _1981_[6:2], _1794_ };
  assign { _2037_[80:26], _1823_, _2037_[24:21], _1515_, _2037_[19:0] } = { _1999_[120], _1109_, _1999_[118:100], _1030_, _1999_[98:76], _1817_, _1999_[74:67], _0574_, _1999_[65:40] } + { _2038_[80:48], _1039_, _2038_[46], _0092_, _2038_[44:43], _0630_, _0407_, _2038_[40:25], _1060_, _2038_[23:11], _2034_[23:15], _2038_[1:0] };
  assign { _1941_[13:1], _0895_ } = { _2039_[13:11], _1417_, _0566_, _1464_, _0581_, _0455_, _0042_, _0518_, _0241_, _1368_, _0795_, _1550_ } + { _1795_, _1014_, _1952_[141], _1621_, _1577_, _1320_, _1952_[137], _0242_, _0109_, _1127_, _0730_, _0318_, _0587_, _0251_ };
  assign { _2001_[111], _1323_, _2001_[109], _1309_, _1081_, _2001_[106:103], _1351_, _2001_[101:99], _1353_, _2001_[97], _1359_ } = { _2014_[14:10], _1988_[54:51], _0291_, _1988_[49], _1383_, _1988_[47:46], _1697_, _0206_ } + in_data[1761:1746];
  assign { _1037_, _1567_ } = { _1966_[32], _0174_ } + { _0299_, _0223_ };
  assign { _1951_[169:159], _1255_, _1951_[157:151], _1276_, _1951_[149:144], _1042_, _1951_[142:139], _0124_, _0929_, _1951_[136:134] } = { _1556_, _0114_, _0319_, _2041_[32:31], _1755_, _2041_[29:24], _0733_, _0915_, _0316_, _0189_, _0194_, _2001_[111], _1323_, _2001_[109], _1309_, _1081_, _2001_[106:103], _1351_, _2001_[101:99], _1353_, _2001_[97], _1359_, _0152_, _1000_, _0356_ } + { in_data[1342:1333], _0043_, _0275_, _0043_, _0082_, _0317_, _2040_[20:11], _0618_, _1485_, _2040_[8], _1488_, _2040_[6:3], _0096_, _0690_, _0068_ };
  assign { _2042_[12:1], _1532_ } = { _2043_[12:2], _0605_, _1009_ } + { _2036_[14], _0509_, _0236_, _2036_[11:3], _1715_ };
  assign { _1431_, _1959_[4:3], _1145_ } = { _0299_, _0324_, _0243_, _0152_ } + { _1225_, _1141_, _0622_, _1986_[1] };
  assign { _2044_[8:6], _0668_, _2044_[4:1], _1461_ } = { _1368_, _0335_, _0646_, _0232_, _0915_, _0905_, _0134_, _0166_, _1352_ } + { _2045_[8:5], _2012_[43:40], _0524_ };
  assign { _1639_, _1900_[46:37], _0767_, _1900_[35:29], _0230_, _1833_, _1900_[26] } = { _1951_[156:151], _1276_, _1951_[149:144], _1042_, _1951_[142:139], _0124_, _0929_, _1951_[136:135] } + { _2038_[27:25], _1060_, _2038_[23:21], _0116_, _0354_, _0522_, _0187_, _0249_, _0217_, _0242_, _0193_, _2046_[6], _1756_, _2046_[4], _1094_, _2046_[2:0] };
  assign { _2047_[83:80], _1445_, _2047_[78:58], _0850_, _2047_[56:14], _1617_, _2047_[12:5], _0679_, _2047_[3:2], _0954_, _2047_[0] } = { _2049_[83:72], _1121_, _2049_[70:69], _2030_[66:46], _0705_, _2030_[44:42], _1598_, _2030_[40:16], _1685_, _2030_[14:0], _0995_, _0082_ } + { _1969_[34:29], _0985_, _1969_[27:15], _0383_, _0186_, _1127_, _0133_, _1994_[9:6], _0840_, _1994_[4:3], _0597_, _2048_[51:50], _1423_, _2048_[48:47], _2005_[10:8], _1327_, _2005_[6:4], _2048_[39:38], _1150_, _2048_[36], _1010_, _2048_[34:17], _0192_, _2023_[13:12], _1469_, _1408_, _2023_[9:7], _0327_, _2023_[5:0], _0425_, _0091_ };
  assign { _2050_[9:5], _1164_, _2050_[3:2], _1296_, _2050_[0] } = { _2051_[9], _1056_, _0121_, _0043_, _0642_, _0161_, _1360_, _0135_, _0146_, _0144_ } + { _1951_[155:151], _1276_, _1951_[149:146] };
  assign { _2052_[40:31], _0252_, _0331_, _2052_[28:17], _0777_, _2052_[15:0] } = { _2054_[40:39], _2039_[13:11], _1417_, _2054_[34:31], _1683_, _2054_[29:19], _1538_, _2054_[17:16], _1029_, _2054_[14:9], _1337_, _2054_[7:2], _1633_, _0156_ } + { _2053_[40:28], _1667_, _2053_[26:21], _1695_, _2053_[19:15], _1185_, _2053_[13:11], _0129_, _0141_, _0152_, _0254_, _1044_, _1066_, _0116_, _0058_, _0071_, _0161_, _0340_ };
  assign { _1415_, _2055_[2:0] } = { _2056_[3:1], _0510_ } + { _1976_[50:49], _0106_, _0191_ };
  assign { _1484_, _1770_, _1935_[47] } = { _2057_[2:1], _1023_ } + in_data[2017:2015];
  assign { _2058_[95:92], _1288_, _2058_[90:60], _1427_, _2058_[58:0] } = { _2033_[20:6], _0196_, _0325_, _2023_[13:12], _1469_, _1408_, _2023_[9:7], _0327_, _2023_[5:0], _0512_, _0023_, _0607_, _1625_, _0627_, _0099_, _2060_[58:51], _0862_, _2060_[49], _2057_[2:1], _2060_[46], _1719_, _2060_[44:40], _1393_, _1136_, _0306_, _0174_, _0657_, _1464_, _0359_, _0019_, _1368_, _1013_, _1266_, _0769_, _0997_, _0979_, _2001_[111], _1323_, _2001_[109], _1309_, _1081_, _2001_[106:103], _1351_, _2001_[101:99], _1353_, _2001_[97], _1359_, _0068_, _0671_, _1589_, _0191_, _1170_, _0003_, _1072_, _0438_, _1625_, _0290_ } + { _2059_[95:89], _0992_, _2059_[87:76], _0547_, _2059_[74:71], _1282_, _2059_[69:67], _1608_, _2059_[65:55], _0822_, _2059_[53:44], _1632_, _2059_[42:32], _1474_, _2059_[30:23], _1330_, _2059_[21:18], _1382_, _2059_[16:6], _1249_, _2059_[4:2], _0697_, _0192_ };
  assign { _2061_[10:4], _1554_, _2061_[2:0] } = { _1971_[22:19], _0922_, _1971_[17:13], _1525_ } + { _2042_[8:1], _0178_, _0924_, _0042_ };
  assign _1942_[86:58] = { _2000_[41:35], _1747_, _2000_[33:31], _1307_, _2000_[29:28], _0303_, _0205_, _0939_, _0654_, _0102_, _0227_, _0144_, _0283_, _1345_, _1358_, _0135_, _0163_, _0278_, _0678_, _0180_ } + { _1982_[7:6], _1287_, _2002_[6:1], _0241_, _0214_, _0243_, _0325_, _0157_, _0206_, _0012_, _0656_, _0332_, _0408_, _1311_, _0287_, _0165_, out_data[416], _0164_, _0018_, _0608_, _1225_, _0228_, _0043_ };
  assign { _2062_[43:28], _0538_, _2062_[26:21], _1849_, _2062_[19:18], _1644_, _2062_[16:6], _1642_, _2062_[4:0] } = { _1890_[11], _0350_, _0228_, _0177_, _0490_, _0552_, _2064_[37], _1350_, _2064_[35:34], _2024_[13:12], _1825_, _2024_[10:2], _2064_[21:14], _1676_, _2064_[12:11], _1049_, _1566_, _2064_[8:7], _0408_, _0343_, _0627_, _1064_, _0572_, _0730_, _0505_ } + { _2063_[43], _1615_, _0147_, _2063_[40:38], _1911_[14:8], _1284_, _0908_, _2063_[28], _0059_, _0179_, _2042_[12:1], _1532_, _0419_, _0217_, _0220_, _0166_, _1343_, _1977_[25:24], _1243_, _1384_, _1669_, _0256_, _0617_, _0129_ };
  assign { _1917_[8:5], _1731_, _1917_[3], _1087_, _1917_[1] } = { _0132_, _0350_, _0609_, _0324_, _0325_, _0133_, _0317_, _0304_ } + { _2057_[1], _2060_[46], _1719_, _2060_[44:43], _0272_, _0454_, _0015_ };
  assign { _2065_[57:40], _1400_, _2065_[38:27], _1430_, _2065_[25:0] } = { _2029_[31:30], _1012_, _2029_[28:19], _1357_, _2029_[17], _1440_, _2029_[15:11], _1115_, _2029_[9:1], _1077_, _0248_, _1684_, _2028_[3], _1326_, _2028_[1], _1415_, _2055_[2:0], _0175_, _1311_, _0046_, _1415_, _2055_[2:0], _1170_, _0092_, _1336_, _0012_, _1147_, _0158_, _0841_, _1015_, _1391_, _0228_ } + { _0540_, _0666_, _0122_, _0250_, _2064_[11], _1049_, _1566_, _2064_[8:7], _0683_, _1991_[55:47], _1193_, _1553_, _1991_[44:43], _2031_[33:31], _1788_, _2031_[29:23], _0514_, _2031_[21:19], _1887_[16], _2031_[17], _1101_, _1814_, _2031_[14:3], _1509_, _1235_, _1072_, _1206_ };
  assign { _2066_[9:6], _1937_, _1736_, _1480_, _2066_[1:0] } = _1968_[44:35] + { _2027_[9], _0042_, _0924_, _1059_, _1393_, _0648_, _1028_, _0726_, _1020_, _0914_ };
  assign { _2068_[32:31], _1058_, _2068_[29:0] } = { _2070_[32:18], _1201_, _2070_[16:11], _1796_, _2070_[9:5], _0165_, _2070_[3:1], _0166_ } + { _2069_[32:23], _1317_, _2069_[21:13], _0202_, _0226_, _0531_, _1680_, _2069_[8], _1458_, _2069_[6:5], _0696_, _1649_, _2069_[2], _0325_, _0922_ };
  assign { _0926_, _0674_, _0610_, _2067_[2:1], _0775_ } = { _1365_, _0104_, _1476_, _1467_, _0277_, _0915_ } + { _0128_, _0103_, _0638_, _0134_, _0317_, _0127_ };
  assign { _1901_[66:63], _1575_, _1901_[61] } = { _2023_[7], _0327_, _2023_[5:2] } + { _1999_[83:82], _0166_, _0615_, _0003_, _0134_ };
  assign { _1936_[47:44], _1612_, _1936_[42], _0418_, _1936_[40] } = { _0024_, _0683_, _0287_, _0274_, _0228_, _0014_, _0306_, _0489_ } + { _1946_[2], _1086_, _0332_, _0953_, _0919_, _0611_, _0989_, _0585_ };
  assign { _2071_[44:37], _1824_, _2071_[35:22], _1900_[86:79], _2071_[13:6], _0427_, _2071_[4:0] } = { _1941_[13:1], _0895_, _1127_, _0058_, _0209_, _1004_, _0408_, _1971_[25:19], _0922_, _1971_[17:13], _1525_, _1971_[11:0] } + { _2072_[44], _1973_[25:24], _0504_, _1597_, _0684_, _1973_[20:19], _1970_[51:42], _1013_, _0662_, _0505_, _0277_, _2040_[20:11], _0618_, _1485_, _2040_[8], _1488_, _2040_[6:3], _1322_, _0661_, _1374_, _1035_, _0175_ };
  assign { _2073_[6:5], _0973_, _2073_[3], _0280_, _2073_[1:0] } = { _2074_[6], _2049_[83:82], _0246_, _0865_, _0354_, out_data[1920] } + { _0692_, _0229_, _0587_, _0503_, _0651_, _0241_, _0905_ };
  assign { _2075_[14:8], _0832_, _2075_[6], _0927_, _2075_[4:0] } = { _1988_[41:40], _1632_, _2027_[10:9], _0889_, _2027_[7:5], _0260_, _2027_[3:1], _1107_, _1038_ } + { _2001_[95:87], _0641_, _0356_, _0289_, _1374_, _0005_, _0016_ };
  assign { _2076_[28:23], _1610_, _2076_[21:0] } = { _1999_[105:100], _1030_, _1999_[98:77] } + { _0364_, _1888_[13], _0036_, _0706_, _1888_[10], _1099_, _0425_, _0110_, _0994_, _0146_, _0578_, _0722_, _0356_, _0194_, _0232_, _0503_, _1144_, _0058_, _0726_, _1027_, _0068_, _0613_, _0652_, _0529_, _0848_, _0368_, _0018_, _0690_, _0746_ };
  assign { _2077_[20], _1403_, _2077_[18:15], _0742_, _2077_[13:10], _0089_, _2077_[8:7], _1227_, _1643_, _1542_, _2077_[3:0] } = { _0581_, _0148_, _0489_, _0221_, _0619_, _0752_, _2042_[12:1], _1532_, _0637_, _0891_ } + { _1975_[74:61], _1786_, _0402_, _1397_, _1569_, _1970_[5], _0681_, _0139_ };
  assign { _2078_[21:16], _0579_, _1173_, _2078_[13:6], _0826_, _2078_[4:0] } = { _2030_[62:51], _0619_, _0408_, _0177_, out_data[1920], _1362_, _1004_, _0024_, _0173_, _0417_, _0657_ } + { _2079_[21:4], _0228_, _0613_, _0732_, _1015_ };
  assign { _2080_[31:23], _0008_, _2080_[21:8], _1707_, _2080_[6:4], _0974_, _2080_[2:0] } = { _2035_[2], _2082_[30:27], _0628_, _2082_[25:24], _1223_, _2082_[22:19], _1355_, _2082_[17:15], _0025_, _0044_, _0149_, _0379_, _0607_, _1936_[47:44], _1612_, _1936_[42], _0418_, _1936_[40], _0619_, _0009_ } + { _1911_[14:8], _1284_, _0908_, _2063_[28], _2081_[21], _1269_, _2081_[19], _1376_, _2081_[17:16], _0127_, _0337_, _0134_, _1633_, _0662_, _0988_, _0091_, _1627_, _0285_, _0999_, _1901_[66:63], _1575_, _1901_[61] };
  assign { _1913_[36:31], _1466_, _1913_[29:25], _0567_, _1701_, _1913_[22:10], _1821_, _1913_[8] } = { _1988_[34:27], _1406_, _0140_, _0220_, _0924_, _1530_, _0588_, _1890_[11], _0350_, _0716_, _1890_[8:6], _0294_, _0228_, _1026_, _0058_, _0307_, _0101_, _0153_, _0261_, _1019_ } + { _2083_[28:7], _0361_, _0716_, _0163_, _0512_, _0681_, _1447_, _0198_ };
  assign { _2084_[9:7], _1906_[4:1], _0744_, _2084_[1], _1420_ } = { _2085_[9], _2074_[6], _2049_[83:78], _0394_, _0650_ } + { _2017_[55:51], _0655_, _0127_, _0453_, _0191_, _0354_ };
  assign { _1935_[79], _1157_, _1935_[77:72], _1953_[24:8], _1428_, _1953_[6], _1776_, _2086_[3:0] } = { _2062_[33:28], _0538_, _2062_[26:21], _1849_, _2062_[19:18], _1644_, _2062_[16:10], _0671_, _0848_, _0099_, _0145_, _0419_, _0014_, _0232_, _0080_ } + { _2087_[31], _1966_[4], _0818_, _1966_[2], _0394_, _0092_, _0401_, _0140_, _1033_, _0228_, _2077_[20], _1403_, _2077_[18:15], _0742_, _2077_[13:10], _0089_, _2077_[8:7], _1227_, _1643_, _1542_, _2077_[3:0], _1689_ };
  assign { _2088_[22:20], _0577_, _2088_[18:0] } = { _1943_[22:5], _0647_, _1943_[3:2], _0018_, _1799_ } + { _2077_[20], _1403_, _2077_[18:15], _0742_, _2077_[13:10], _0089_, _2077_[8:7], _1227_, _1643_, _1542_, _2077_[3:0], _0631_, _1368_ };
  assign { _1716_, _1996_[4], _1365_, _0104_, _1476_, _1467_ } = { _0189_, _0025_, _0250_, _0154_, _0025_, _0189_ } + { _0101_, _0025_, _0241_, _0356_, _0356_, _0025_ };
  assign { _2089_[5:4], _1769_, _2089_[2], _1526_, _0011_ } = { _1900_[45:41], _1405_ } + { _1952_[14:12], _1385_, _1952_[10], _0643_ };
  assign { _2090_[14:11], _1945_[7:5], _1519_, _2090_[6:0] } = { _2092_[14:7], _1548_, _2092_[5], _2064_[11], _1049_, _1566_, _2064_[8:7] } + { _2091_[14:13], _0644_, _2091_[11], _2014_[17:10], _1174_, _0550_, _0924_ };
  assign { _2093_[130:128], _1071_, _2093_[126:77], _1591_, _2093_[75:55], _1899_[53:3], _2093_[3:0] } = { _2095_[130:127], _2007_[8:1], _1441_, _2095_[117:108], _1972_[25:23], _1686_, _0335_, _0076_, _1981_[11:9], _0299_, _0223_, _1981_[6:2], _1794_, _0189_, _0190_, _0694_, _0127_, _2095_[86:40], _1516_, _2095_[38:26], _1352_, _2095_[24], _1661_, _1710_, _2095_[21], _1162_, _1272_, _2095_[18:12], _1585_, _0746_, _0466_, _0338_, _0784_, _0946_, _0703_, _1225_, _0619_, _0907_, _0419_, _0678_ } + { _2094_[130:103], _1291_, _2094_[101:94], _1263_, _2094_[92:69], _0246_, _0332_, _0549_, _1195_, _0179_, _0183_, _0210_, _0303_, _0999_, _0598_, _0702_, _0612_, _0106_, _2094_[55:47], _1732_, _2094_[45], _1283_, _0103_, _2046_[6], _1756_, _2046_[4], _1094_, _2046_[2:0], _0043_, _0191_, _0151_, _1044_, _0704_, _0288_, _1021_, _2094_[28:26], _1779_, _2094_[24], _0691_, _1416_, _1781_, _2094_[20:19], _0545_, _2094_[17:14], _0346_, _2094_[12:6], _1767_, _2094_[4:3], _1645_, _0043_, _1799_ };
  assign _2096_ = { _1984_[41:39], _1714_, _1984_[37:36], _0251_, _1984_[34:26], _1005_, _0057_, _1044_, _0808_, _1468_, _2098_[18:3], _0289_, _0206_, _1392_ } + { _2097_[39:5], _1037_, _1567_, _0299_, _0069_, _0032_ };
  assign { _2099_[9], _1840_, _2099_[7], _1426_, _2099_[5:0] } = { _1987_[40:37], _1402_, _0656_, _0041_, _0356_, _0271_, _0057_ } + { _1357_, _2029_[17], _1440_, _2029_[15], _0709_, _0225_, _0096_, _0708_, _0695_, _1114_ };
  assign { _2100_[165:28], _0508_, _2100_[26:0] } = { _0865_, _1651_, _0134_, _0289_, _0683_, _0681_, _0984_, _1247_, _0221_, _2096_, _0642_, _2102_[115:53], _0399_, _2102_[51:34], _1662_, _2102_[32:13], _2073_[6:5], _0973_, _2073_[3], _0280_, _2073_[1:0], _0521_, _0692_, _0137_, _0681_, _0978_, _0631_ } + { _2101_[165:163], _2045_[8:5], _2012_[43:28], _1625_, _2012_[26:22], _1678_, _1222_, _2012_[19:2], _1613_, _2101_[115:111], _1368_, _0566_, _1951_[123], _1122_, _1951_[121:119], _1609_, _0379_, _0096_, _1395_, _1380_, _0603_, _0152_, _0626_, _0683_, _1392_, _2101_[93:90], _0910_, _2101_[88], _1895_[35:26], _1111_, _1895_[24:20], _1757_, _1895_[18:3], _1634_, _0166_, _0752_, _1655_, _0198_, _0642_, _0438_, _0204_, _2101_[46:40], _1163_, _2101_[38:34], _1216_, _2101_[32:27], _0658_, _1980_[23:6], _1367_, _1980_[4], _1681_, _1980_[2:0], _0518_, _0914_ };
  assign _2103_ = { _0117_, _0710_, _0519_, _0228_, _0450_, _0239_, _1401_ } + { _2104_[6:3], _0648_, _0354_, _1283_ };
  assign { _2000_[123:108], _1361_, _2000_[106:100], _1506_, _2000_[98], _0113_, _2000_[96:92], _0313_, _2000_[90:86], _0737_, _2000_[84:80] } = { _2105_[43:38], _2035_[23:19], _1455_, _1507_, _2035_[16], _1674_, _2035_[14:2], _2082_[30:27], _0628_, _2082_[25:24], _1223_, _2082_[22:19], _1355_, _0265_, _1000_, _0238_ } + { _2025_[43:40], _1785_, _2025_[38:34], _1510_, _2025_[32:27], _0896_, _2025_[25], _1556_, _0114_, _0319_, _2041_[32:31], _0356_, _0250_, _0154_, _0661_, _0152_, _1046_, _0661_, _1283_, _0152_, _0152_, _0134_, _0226_, _0084_, _0084_, _0138_, _0317_, _0356_, _0733_, _0043_, _0277_ };
  assign { _2106_[30:25], _1728_, _2106_[23:22], _0040_, _2106_[20:0] } = { _1995_[14], _0224_, _1995_[12], _1379_, _0041_, _2069_[8], _1458_, _2069_[6:5], _0696_, _1649_, _2069_[2], _0175_, _0176_, _1020_, _1601_, _2107_[14:13], _2092_[14:7], _1548_, _2092_[5], _2107_[2:1], _0368_ } + { _1967_[6:1], _2078_[21:16], _0579_, _1173_, _2078_[13:6], _0826_, _2078_[4:0], _1689_, _1645_, _0904_ };
  assign { _2109_[8:1], _1546_ } = { _2068_[19:17], _0636_, _0718_, _0284_, _0456_, _0631_, _0000_ } + { _2050_[2], _1296_, _2050_[0], _0686_, _0297_, _0351_, _0454_, _0018_, _1132_ };
  assign { _2110_[51:46], _1103_, _2110_[44:0] } = { _1503_, _2111_[50:35], _0661_, _2111_[33:29], _2087_[31], _2111_[27:21], _1200_, _2111_[19:4], _0489_, _0469_, _1702_, _0866_ } + { _2094_[126:103], _1291_, _2094_[101:94], _1263_, _2094_[92:75] };
  assign { _2113_[25:11], out_data[544], _1933_[28:19] } = { _2114_[25:23], _0189_, _0759_, _1976_[19:16], _1335_, _1976_[14], _0172_, _0120_, _1568_, _1976_[10:9], _0604_, _1976_[7], _0945_, _1976_[5], _0602_, _1976_[3:0], _0857_ } + { _2058_[39:22], _1051_, _0752_, _0245_, _0652_, _0290_, _0253_, _0716_, _0234_ };
  assign { _2115_[14:8], _1479_, _1924_[7], _0847_, _2115_[4:2], _0869_, _2115_[0] } = { _2000_[118:108], _1361_, _2000_[106], _0284_, _0740_ } + { _1952_[42], _0803_, _1952_[40:33], _0202_, _0977_, _0307_, _0594_, _0146_ };
  assign { _2116_[8], _1499_, _2116_[6:5], _1448_, _2116_[3], _1523_, _2116_[1:0] } = { _2117_[8:6], _0432_, _2117_[4:1], _0607_ } + { _1968_[25:19], _0121_, _1363_ };
  assign _2118_ = { _1157_, _1935_[77:72], _1953_[24:8], _1428_, _1953_[6], _1776_, _0482_, _1761_, _1590_, _1929_[4:3], _1073_, _1627_, _1026_, _1409_, _2106_[30:25], _1728_, _2106_[23:22], _0040_, _2106_[20:0], _2120_[32:30], _1762_, _2120_[28:16], _0793_, _1425_, _1900_[72:70], _0389_, _1900_[68:66], _0833_, _1305_, _1900_[63], _0159_, _0466_, _0299_, _0924_ } + { _2038_[39:31], _0323_, _2080_[31:23], _0008_, _2080_[21:8], _1707_, _2080_[6:4], _0974_, _2080_[2:0], _0781_, _0559_, _0068_, _0059_, _1551_, _0228_, _0000_, _0857_, _1421_, _0265_, _0887_, _0113_, _0014_, _1704_, _0161_, _0671_, _0590_, _0217_, _0216_, _0605_, _2119_[37:30], _1450_, _1638_, _2119_[27:26], _1502_, _2119_[24:20], _0828_, _2051_[9], _2119_[17], _1106_, _2119_[15:14], _1171_, _2119_[12:3], _0030_, _0272_, _0631_ };
  assign { _2122_[22:9], _1949_[9:5], _1273_, _2122_[2:0] } = { _2123_[22:1], _0129_ } + { _2100_[84:68], _0264_, _1425_, _0662_, _0149_, _0944_, _0383_ };
  assign { _2124_[14:9], _1452_, _1964_[75:74], _1647_, _1964_[72:68] } = { _2065_[51:40], _1400_, _1004_, _0014_ } + { _2119_[20], _0828_, _2051_[9], _2119_[17], _1106_, _2119_[15:14], _1171_, _2119_[12:8], _0736_, _0080_ };
  assign { _2112_[97:95], _1803_, _2112_[93:81], _2095_[130:127], _2007_[8:1], _1441_, _2095_[117:108], _1972_[25:22], _1687_, _1972_[20:11], _2112_[42:28], _1666_, _2112_[26:15], _0262_, _2112_[13:12], _1604_, _2112_[10:6], _0410_, _2112_[4:0] } = { in_data[2137:2084], _2121_[43:39], _0864_, _1346_, _2121_[36:35], _1600_, _2121_[33:28], _0653_, _2121_[26:22], _2031_[66], _0328_, _2031_[64], _0007_, _1699_, _2031_[61:55], _1806_, _2031_[53], _0206_, _2031_[51], _1800_, _2031_[49:47], _2121_[1:0] } + { in_data[1737:1660], _0189_, _0101_, _0356_, _0189_, _0200_, _0241_, _0356_, _0025_, _1716_, _1996_[4], _1365_, _0104_, _1476_, _1467_, _1716_, _1996_[4], _1365_, _0104_, _1476_, _1467_ };
  assign { _2125_[48:44], _0845_, _2125_[42:13], _1277_, _2125_[11:0] } = { _1699_, _2031_[61:59], _2126_[44:43], _2101_[93:90], _0910_, _2101_[88], _1895_[35:26], _1111_, _1895_[24:20], _1757_, _1895_[18:3], _1027_, _0010_, _1554_, _1689_ } + { _2032_[22:19], _0304_, _1392_, _1063_, _1093_, _0032_, _1943_[81:75], _1082_, _1943_[73:68], _1504_, _1943_[66:64], _1724_, _1943_[62:60], _0922_, _2023_[13:12], _1469_, _1408_, _2023_[9:7], _0327_, _2023_[5:0], _1374_, _0401_, _1425_ };
  assign { _2127_[6:2], _1881_, _2127_[0] } = { _1943_[81:78], _1348_, _0238_, _1551_ } + { _2015_[7:2], _1369_ };
  assign { _1942_[16:15], _1279_, _1942_[13:10], _1619_, _1942_[8:4] } = { _2047_[56:47], _0463_, _0670_, _0897_ } + { _2080_[19:10], _0005_, _0153_, _0227_ };
  assign { _2128_[16:2], _0782_, _2128_[0] } = _2129_ + { _2110_[51:46], _1103_, _2110_[44:37], _1179_, _0227_ };
  assign { _1838_, _2130_[5:4], _1492_, _1119_, _0952_, _2130_[0] } = { _0295_, _1208_, _0779_, _0764_, _0215_, _0279_, _0071_ } + { _1164_, _2050_[3:2], _0301_, _0144_, _0261_, _1421_ };
  assign _2131_ = { _0058_, _1818_ } + { _2132_[1], _0282_ };
  assign { _2133_[6:1], _1727_ } = { _1995_[15:14], _0224_, _1995_[12:9] } + { _2134_[6], _0003_, _2134_[4:3], _0530_, _0018_, _0254_ };
  assign _2135_ = { _1849_, _2062_[19:18], _0634_, _0102_, _0034_, _0621_, _0488_ } + { _0140_, _1518_, _0204_, _0356_, _0726_, _1589_, _0530_, _0105_ };
  assign _2136_ = { _1999_[103:101], _0024_, _0745_, _1528_, _0649_, _0025_, _1342_ } + { _2101_[40], _1163_, _2101_[38:34], _1216_, _2101_[32] };
  assign _2137_ = _2052_[6:4] + { _1037_, _1567_, _0242_ };
  assign { _2138_[72:36], _1844_, _2138_[34:0] } = { _2013_[15:10], _1857_, _2013_[8:7], _1829_, _1040_, _2013_[4], _0379_, _0097_, _0009_, _0891_, _0096_, _0633_, _0162_, _1959_[7], _1202_, _1980_[23:6], _1367_, _1980_[4], _1681_, _1980_[2:0], _2139_[26:1], _0454_, _0751_ } + { _1901_[66:63], _1575_, _1901_[61], _2139_[66:60], _1705_, _2139_[58:55], _1743_, _0943_, _2139_[52:51], _0345_, _2139_[49], _1748_, _2139_[47:45], _1837_, _2139_[43], _1256_, _2139_[41:40], _0337_, _1251_, _0590_, _0348_, _2139_[35:32], _1354_, _1054_, _2139_[29:1], _0277_ };
  assign { _1951_[29:6], _0382_, _1951_[4:2] } = { _2066_[8:6], _1937_, _1736_, _1480_, _2066_[1:0], _0489_, _1088_, _2001_[111], _1323_, _2001_[109], _1309_, _1081_, _2001_[106:103], _1351_, _2001_[101:99], _1353_, _2001_[97], _1359_, _0746_ } + { _2058_[71:66], _0702_, _1171_, _0190_, _0190_, _0640_, _0454_, _0015_, _0615_, _1095_, _0285_, _1089_, _0675_, _1421_, _1147_, _0707_, _1609_, _0259_, _1424_, _0081_, _1340_, _0018_, _0675_ };
  assign { _1956_[30:24], _1618_, _1956_[22], _2140_[13:0] } = { _2060_[58:51], _0862_, _1964_[52], _1795_, _1964_[50:48], _1016_, _1964_[46:45], _0492_, _1964_[43], _1706_, _0226_, _0700_, _1028_ } + { _2141_[22:19], _1901_[15:14], _0760_, _1901_[12:10], _0879_, _1901_[8:5], _1078_, _1901_[3], _0660_, _0311_, _1651_, _0057_, _0530_, _1017_ };
  assign { _2147_[5], _1869_, _2147_[3:0] } = _2146_[13:8] + _2058_[65:60];
  assign { _2148_[60:50], _1851_, _2148_[48:39], _0880_, _2148_[37:30], _1934_[5:4], _2148_[27:7], _1578_, _2148_[5:0] } = { _2143_[36:3], _2150_[26:0] } + { _2149_[60:20], _1063_, _0228_, _0680_, _0305_, _1064_, _0228_, _2149_[13:8], _1152_, _2149_[6], _0258_, _0297_, _1360_, _0132_, _0685_, _1363_ };
  assign { _1891_[12:5], _2144_[55], _1250_, _2072_[44], _1973_[25:24], _0504_, _1597_, _0684_, _1973_[20:19], _1970_[51:20], _1253_, _1970_[18:16], _1210_, _1682_, _1970_[13:11], _2144_[4:0] } = { _2112_[87:81], _2095_[130:127], _2007_[8:1], _1441_, _2095_[117:108], _1972_[25:22], _1687_, _1972_[20:11], _2112_[42:28], _1666_, _2112_[26:25], _0058_ } + { _2112_[85:81], _2095_[130:127], _2007_[8:1], _1441_, _2095_[117:108], _1972_[25:22], _1687_, _1972_[20:11], _2112_[42:28], _1666_, _2112_[26:22] };
  assign _2152_ = { _2029_[1], _0189_, _0663_, _1818_ } + { _2126_[44:43], _0710_, _0359_ };
  assign { _2000_[20:19], _0564_, _2000_[17:14], _0925_, _1939_[12:8], _0501_, _1939_[6], _1306_, _2000_[4:3], _1632_, _1373_, _2000_[0] } = { _2041_[26:24], _0233_, _0499_, _2114_[25:24], _0043_, _0219_, _0125_, _1235_, _0043_, _0191_, _0134_, _0907_, _0608_, _1206_, _0058_, _0317_, _1211_, _1393_ } + { _1972_[19:16], _0097_, _0121_, _0401_, _1203_, _0356_, _0152_, _0106_, _0241_, _0690_, _1235_, _1046_, _0926_, _0674_, _0610_, _2067_[2:1], _0775_ };
  assign { _2153_[39:24], _1508_, _2153_[22:0] } = { _0563_, _0620_, _0993_, _0403_, _1935_[79], _1157_, _1935_[77:72], _1953_[24:8], _1428_, _1953_[6], _1776_, _2086_[3:0], _1329_, _1000_, _0612_, _0265_ } + { _2154_[39:35], _1080_, _2154_[33:32], _1338_, _0851_, _0242_, _0540_, _0318_, _0417_, _2044_[8:6], _0668_, _2044_[4:1], _1461_, _0905_, _0323_, _0076_, _1941_[13:1], _0895_ };
  assign { _2155_[11:2], _1871_, _2155_[0] } = { _2025_[31], _0081_, _1340_, _1019_, _0250_, _0995_, _0241_, _0466_, _0321_, _1043_, _0251_, _0116_ } + _2068_[29:18];
  assign _2156_ = { _2017_[64:61], _1364_, _2017_[59:37], _1410_, _2017_[35:33], _0414_, _2017_[31:14], _1442_, _2017_[12:6], _1810_, _0123_, _1932_[6], _0595_, _0311_, _0335_, _0295_, _0915_, _1912_[29:15], _1592_, _1912_[13:10], _0188_, _1912_[8:2], _0967_, _0134_, _0723_, _0155_, _1974_[0], _1174_, _0450_, _0883_ } + { _2094_[122:103], _1291_, _2094_[101:97], _0023_, _1977_[25:24], _1243_, _1384_, _1669_, _0256_, _0811_, _0145_, _0453_, _0106_, _2136_, _0477_, _0144_, _0986_, _1908_[14:13], _1564_, _1908_[11:10], _0535_, _1908_[8:7], _0979_, _2108_[80:78], _1791_, _2108_[76], _2053_[40:28], _1667_, _2053_[26:21], _1695_, _2053_[19:15], _1185_, _2053_[13:11], _2108_[45:43], _0071_, _0153_, _0102_, _0724_, _0566_, out_data[1600], _1371_ };
  assign _2157_ = { _2148_[57:50], _1851_, _2148_[48:39], _0880_, _2148_[37:30], _0887_, _1105_, _0116_, _0003_, _0284_, _0642_, _1007_, _0000_, _1457_, _0071_, _0354_ } + { _1376_, _2119_[37:30], _1450_, _1638_, _2119_[27:26], _1502_, _2119_[24:20], _0828_, _2051_[9], _2119_[17], _1106_, _2119_[15:14], _1171_, _2119_[12:3], _1812_, _0018_, _0458_ };
  assign { _0633_, _0162_, _1959_[7], _1202_ } = { _0350_, _0716_, _0191_, _0383_ } + { _0926_, _0674_, _0610_, _2067_[2] };
  assign { _1539_, _1935_[26:25] } = { _0279_, _0175_, _0287_ } + { _1366_, _0768_, _0128_ };
  assign { _2158_[50:48], _1300_, _2158_[46:40], _1563_, _2158_[38:34], _1489_, _2158_[32:0] } = { _2160_[50:24], _0749_, _0590_, _1901_[66:63], _1575_, _1901_[61], _0855_, _1459_, _0058_, _0298_, _1936_[47:44], _1612_, _1936_[42], _0418_, _1936_[40], _1121_, _0366_, _0548_, _0649_ } + { _2159_[50:48], _1907_[55:25], _1535_, _1907_[23:16], _2159_[7:2], _1842_, _2159_[0] };
  assign { _2162_[42:18], _0874_, _2162_[16], _1766_, _2162_[14:9], _1155_, _2162_[7:0] } = { _2030_[50:46], _0705_, _2030_[44:42], _1598_, _2030_[40:16], _1685_, _2030_[14:8] } + { _2163_[42:25], _0228_, _1228_, _0748_, _1655_, _1051_, _0703_, _1088_, _1348_, _0566_, _0358_, _0936_, _0221_, _1090_, _0323_, _1951_[123], _1122_, _1951_[121:119], _1609_, _0267_, _0899_, _0279_, _0034_, _0988_ };
  assign { _2164_[29:24], _0601_, _2164_[22:20], _1997_, _2164_[16:12], _2154_[39:35], _1080_, _2154_[33:32], _1338_, _2164_[2:0] } = { _2000_[123:108], _1361_, _2000_[106:100], _0152_, _0518_, _0237_, _1551_, _0097_, _0354_ } + { _1393_, _0232_, _0661_, _0128_, _0993_, _0403_, _0993_, _0403_, _0586_, _0219_, _0058_, _2040_[20:11], _0618_, _1485_, _2040_[8], _1488_, _2040_[6:3], _0661_ };
  assign { _1887_[14], _0852_, _1887_[12] } = { _0047_, _0027_, _0213_ } + { _1049_, _0013_, _0642_ };
  assign { _2167_[6], _1524_, _2167_[4:0] } = { _0380_, _0728_, _0825_, _0694_, _0300_, _0678_, _0041_ } + _2032_[21:15];
  assign { _1991_[55:47], _1193_, _1553_, _1991_[44:43], _2031_[33:31], _1788_, _2031_[29:23], _0514_, _2031_[21:19], _1887_[16], _2031_[17], _1101_, _1814_, _2031_[14:3], _1509_ } = { _0219_, _0189_, _0022_, _1677_, _0409_, _1804_, _1386_, _2002_[27:26], _1381_, _1520_, _1982_[21:16], _1534_, _1982_[14:6], _1287_, _2002_[6:0], _0306_, _1235_, _0306_, _0116_, _0146_, _0633_, _0162_, _1959_[7], _1202_, _0025_ } + { _1952_[191:184], _1389_, _1952_[182:177], _0344_, _1952_[175:165], _0311_, _2001_[111], _1323_, _2001_[109], _1309_, _1081_, _2001_[106:103], _1351_, _2001_[101:99], _1353_, _2001_[97], _1359_, _0272_ };
  assign { _2168_[169:166], _1521_, _2168_[164:111], _1989_[54:33], _1344_, _1989_[31:5], _1792_, _1989_[3:2], _1992_[8], _2168_[56:0] } = { _2000_[122:108], _1361_, _2000_[106:100], _1506_, _2000_[98], _0113_, _2000_[96:92], _0313_, _2000_[90:86], _0737_, _2000_[84:83], _0237_, _1206_, _0573_, _1046_, _0084_, _0270_, _0464_, _0638_, _0272_, _0356_, _0232_, _1283_, _0071_, _2164_[29:24], _0601_, _2164_[22:20], _1997_, _2164_[16:12], _2154_[39:35], _1080_, _2154_[33:32], _1338_, _2164_[2:0], _0194_, _0317_, _2170_[84:70], _2070_[32:18], _1201_, _2070_[16:11], _1796_, _2070_[9:5], _0165_, _2070_[3:1], _2170_[37:31], _1008_, _2170_[29:26], _1332_, _2170_[24:9], _0169_, _2170_[7:4], _1203_, _0354_, _0232_, _0241_ } + { _1972_[13:11], _2112_[42:28], _1666_, _2112_[26:15], _0262_, _2112_[13:12], _1604_, _2112_[10:6], _0410_, _2112_[4:1], _1203_, _0189_, _0228_, _0189_, _1153_, _1893_[10:7], _1034_, _1893_[5:4], _1374_, _1787_, _0126_, _1328_, _0287_, _0238_, _0134_, _0304_, _0205_, _0096_, _0200_, _2169_[101], _2105_[43:38], _2035_[23:19], _1455_, _1507_, _2035_[16], _1674_, _2035_[14:2], _2082_[30:27], _0628_, _2082_[25:24], _1223_, _2082_[22:19], _1355_, _2082_[17:15], _2169_[56:55], _0451_, _2169_[53:45], _1793_, _2169_[43:40], _1324_, _2169_[38:35], _2000_[59:50], _1570_, _2000_[48:46], _1314_, _1419_, _0391_, _2000_[42:35], _1747_, _2000_[33:31], _1307_, _2000_[29:27], _1318_, _0106_ };
  assign _2171_ = { _1912_[19], _0168_, _1088_ } + { _1985_[3], _1841_, _0849_ };
  assign _2172_ = { _2071_[44:37], _1824_, _2071_[35:28], _0046_, _0700_, _1843_, _1733_, _0096_, _0282_, _0286_ } + { _2173_[23:21], _1460_, _2173_[19:3], _0163_, _1443_, _1471_ };
  assign { _2174_[9], _0444_, _1572_, _1653_, _2174_[5:2], _0969_, _2174_[0] } = { _0487_, _0324_, _0736_, _0549_, _2137_, _0071_, _0995_, _0342_ } + { _1079_, _0726_, _0243_, _0752_, _0058_, _0353_, _1356_, _1472_, _0348_, _0149_ };
  assign { _2175_[12:7], _1252_, _2175_[5:4], _0839_, _0836_, _2175_[1:0] } = { _2143_[62:53], _0600_, _0553_, _0987_ } + { _2029_[20:19], _1357_, _0338_, _1810_, _0123_, _1932_[6], _0595_, _0079_, _0116_, _0033_, _0866_, _1274_ };
  assign _2179_ = { _1940_[22:20], _1901_[86:85], _0949_, _1439_ } + _2180_;
  assign { _2182_[102:77], _1925_[30:7], _2182_[52:43], _0584_, _2182_[41:26], _0976_, _2182_[24:0] } = { _2183_[102:50], _1349_, _2183_[48:29], _2079_[21:16], _0571_, _1977_[25:24], _1243_, _1384_, _1669_, _0256_, _0041_, _1720_, _0656_, _2183_[12:9], _0906_, _2183_[7:3], _0044_, _0888_, _0367_ } + { _2093_[111:77], _1591_, _2093_[75:55], _1899_[53:13], _0179_, _1729_, _1133_, _1847_, _0808_ };
  assign { _2184_[13], _1630_, _2184_[11:6], _1740_, _2184_[4:0] } = { _2038_[35:34], _0119_, _1900_[72:70], _0389_, _1900_[68:66], _0833_, _1305_, _1900_[63], _1501_ } + { _2001_[88:86], _0998_, _2001_[84:78], _1031_, _0550_, _1381_ };
  assign { _1964_[32:31], _1156_, _1964_[29:27] } = { _1539_, _1935_[26:25], _0326_, _1290_, _0637_ } + _2093_[126:121];
  assign { _2187_[24:23], _1941_[37:24], _2187_[8:4], _1745_, _2187_[2:0] } = { _2185_[37:32], _2176_, _1475_, _2185_[22:14], _1299_ } + { _2188_[24:19], _0459_, _2188_[17:5], _0352_, _1691_, _0176_, _1422_, _0796_ };
  assign { _1966_[44:42], _1236_ } = { _0565_, _0571_, _0680_, _0231_ } + { _0629_, _1726_, _0279_, _0795_ };
  assign { _2189_[78:72], _1923_[7:5], _2189_[68:44], _1641_, _2189_[42:37], _1159_, _2189_[35:34], _1588_, _2189_[32:0] } = { _1144_, _0289_, _1579_, _1573_, _2190_[74], _0071_, _1478_, out_data[1184], _0560_, _1129_, _0565_, _0599_, _0206_, _0754_, _0529_, _1009_, _0043_, _1102_, _0633_, _0162_, _1959_[7], _1202_, _2116_[8], _1499_, _2116_[6:5], _1448_, _2116_[3], _1523_, _2116_[1:0], _0325_, _1425_, _1286_, _0511_, _0872_, _2174_[9], _0444_, _1572_, _1653_, _2174_[5:2], _0969_, _2174_[0], _0343_, _0285_, _1614_, _0695_, _0019_, _1348_, _2077_[20], _1403_, _2077_[18:15], _0742_, _2077_[13:10], _0089_, _2077_[8:7], _1227_, _1643_, _1542_, _2077_[3:0], _0893_, _0420_, _1235_, _0157_, _0358_, _0654_ } + { _2182_[48:43], _0584_, _2182_[41:26], _0976_, _2182_[24:2], _0144_, _0034_, _0813_, _0774_, _0718_, _0342_, _1206_, _1614_, _0310_, _1725_, _1298_, _0797_, _0751_, _0704_, _0562_, _1138_, _1465_, _0801_, _1161_, _0178_, _0286_, _1348_, _0222_, _0272_, _0452_, _1471_, _1512_, _0228_, _0031_, _1438_, _0563_, _1834_ };
  assign { _2191_[9:7], _1914_[46:40] } = { _2176_[5], _0354_, _0239_, _1453_, _0065_, _0780_, _0823_, _1497_, _0371_, _0307_ } + { _2136_[6:1], _0511_, _0424_, _0885_, _0016_ };
  assign { _2192_[37:14], _1944_[35], _2192_[12:0] } = { _2012_[36:28], _1625_, _2012_[26:22], _1678_, _1222_, _2012_[19:2], _1613_, _2101_[115:114] } + { _2100_[34:28], _0508_, _2100_[26:4], _0942_, _0310_, _1235_, _0576_, _0187_, _0339_, _1393_ };
  assign _1894_[18:3] = { _2150_[20:7], _0815_, _0014_ } + { _1982_[18:16], _1534_, _1982_[14:6], _1287_, _0221_, _0405_ };
  assign _2193_ = { _1967_[21:15], _1668_ } + { _0594_, _0756_, _1345_, _0330_, _1464_, _1739_, _1205_, _0059_ };
  assign { _0482_, _1761_, _1590_, _1929_[4:3] } = { _0518_, _0134_, _0311_, _0039_, _0317_ } + { _0250_, _0464_, _0103_, _0150_, _0227_ };
  assign { _1962_[11:5], _1261_, _1962_[3:1] } = { _2195_[10:6], _0412_, _1827_, _1625_, _1610_, _0649_, _0047_ } + { _0726_, _2194_[9], _2134_[6], _0003_, _2134_[4:3], _2194_[4], _0503_, _2165_[11], _1187_, _0004_ };
  assign { _2196_[154:61], _1861_, _2196_[59:0] } = { _2045_[8:5], _2012_[43:28], _1625_, _2012_[26:22], _1678_, _1222_, _2012_[19:9], _1017_, _1172_, _2075_[14:8], _0832_, _2075_[6], _0927_, _2075_[4:0], _2188_[24:19], _0459_, _2188_[17:5], _2187_[24:23], _1941_[37:24], _2187_[8:4], _1745_, _2187_[2:0], _0872_, _0609_, _0733_, _0027_, _0739_, _0700_, _0953_, _0405_, _1411_, _1258_, _0751_, _1134_, _1914_[10], _1529_, _1471_, _1304_, _0809_, _0894_, _0812_, _0267_, _0657_, _0157_, _0587_, _1625_, _0829_, _0824_, _2139_[26:1], _0978_, _0058_ } + { _1971_[24:19], _0922_, _1971_[17:13], _1525_, _1971_[11:3], _0228_, _0285_, _0179_, _0317_, _0631_, _0157_, _1554_, _1468_, _2098_[18:3], _1208_, _1174_, _0704_, _1828_, _0701_, _0298_, _0817_, _0609_, _1017_, _0848_, _0012_, _0009_, _0756_, _0193_, _0217_, _0014_, _0627_, _2197_[91:90], _0877_, _2197_[88:82], _0271_, _0032_, _1481_, _1835_, _2197_[77:26], _0467_, _0337_, _1170_, _1561_, _1456_, _1447_, _1554_, _0669_, _1374_, _0237_, _2152_, _0812_, _1203_, _0368_, _0103_, _0478_, _0027_, _0115_, _0343_, _1585_, _0987_, _1552_, _0709_ };
  assign { _2198_[47:6], _1545_, _2198_[4:0] } = { _2200_[47:42], _1855_, _0923_, _2200_[39:20], _0202_, _1394_, _1046_, _1270_, _0807_, _1154_, _0609_, _2127_[6:2], _1881_, _2127_[0], _0217_, _0670_, _1615_, _0381_, _0347_, _0799_ } + { _2183_[78:59], _2199_[27:21], _0996_, _2199_[19:16], _2010_[3:1], _0240_, _0844_, _1713_, _1433_, _0251_, _2193_ };
  assign { _2202_[4], _1184_, _1773_, _2202_[1], _1774_ } = { _2109_[8:5], _0105_ } + { _0027_, _0873_, _0368_, _0071_, _0238_ };
  assign { _1671_, _2203_[16:10], _1571_, _2203_[8], _1938_[8:5], _0131_, _2203_[2:0] } = { _0113_, _2000_[96:92], _0313_, _2000_[90:86], _0586_, _1786_, _0402_, _1397_, _1569_, _1970_[5] } + { _1982_[7:6], _1287_, _2002_[6:0], _1527_, _0084_, _1786_, _0402_, _1397_, _1569_, _1970_[5], _0311_ };
  assign { _1976_[19:16], _1335_, _1976_[14], _0172_, _0120_, _1568_, _1976_[10:9], _0604_, _1976_[7], _0945_, _1976_[5], _0602_, _1976_[3:0] } = { _2205_[19:18], _0726_, _2194_[9], _2134_[6], _0003_, _2134_[4:3], _2194_[4], _1091_, _2205_[9:3], _1693_, _2205_[1:0] } + { _1615_, _0147_, _2063_[40:38], _1911_[14], _1964_[67], _0364_, _1888_[13], _0036_, _0706_, _1888_[10:5], _0673_, _1964_[55], _1679_ };
  assign _1901_[57:39] = { _1964_[21:10], _1433_, _0733_, _1033_, _0672_, _0134_, _1038_, _1422_ } + { _2175_[12:7], _1252_, _2175_[5:4], _0839_, _0836_, _0377_, _0025_, _0015_, _0779_, _0300_, _0076_, _0454_, _1181_ };
  assign { _2206_[11:7], _0981_, _2206_[5:0] } = { _1909_[39:35], _0254_, _1909_[33:29], _0317_ } + { _0194_, _0222_, _0812_, _1698_, _0225_, _0299_, _2147_[5], _1869_, _2147_[3:0] };
  assign _2207_ = { _1894_[9:7], _0860_, _0277_ } + { _0598_, _2131_, _0393_, _0948_ };
  assign { _2208_[3:1], _1281_ } = { _2179_[2:1], _0308_, _0940_ } + { _1967_[2:0], _0924_ };
  assign { _2210_[13:4], _1875_, _2210_[2:0] } = { _1668_, _1967_[13:10], _1321_, _0473_, _1967_[7], _1204_, _0057_, _1075_, _0641_, _0825_, _0246_ } + { _2211_[13:7], _1541_, _2211_[5:3], _0146_, _1121_, _0687_ };
  assign { _2032_[31:26], _1826_, _2032_[24:13], _0606_, _2032_[11:10], _1754_, _2032_[8:1] } = { _2121_[25:22], _2031_[66], _0328_, _2031_[64], _0007_, _1699_, _2031_[61:55], _1806_, _2031_[53], _0189_, _0482_, _1761_, _1590_, _1929_[4:3], _0633_, _0162_, _1959_[7], _1202_, _0317_, _0221_, _0315_ } + { _0223_, _1981_[6:4], _0134_, _0752_, _0633_, _0162_, _1959_[7], _1202_, _0661_, _0152_, _0857_, _0752_, _0194_, _1283_, _0071_, _0197_, _0518_, _0265_, _0918_, _0219_, _0125_, _0272_, _1170_, _1206_, _0084_, _0290_, _1362_, _1203_, _0603_ };
  assign _1893_[37:14] = { _1490_, _2214_[22], _0034_, _0238_, _2139_[66:60], _1705_, _2139_[58:55], _1743_, _0943_, _2139_[52:51], _0507_, _1139_, _1072_, _1551_ } + { _2213_[23:18], _0208_, _1114_, _1270_, _0192_, _0159_, _1636_, _2117_[8:6], _0432_, _2117_[4:1], _2213_[3], _0347_, _0421_, _1135_ };
  assign { _1947_[11:6], _1267_, _1947_[4:3], _1646_ } = { _2107_[13], _2092_[14:13], _1737_, _1513_, _1454_, _1868_, _1841_, _0433_, _1733_ } + { _2116_[8], _1499_, _2116_[6:5], _1448_, _2116_[3], _1523_, _2116_[1:0], _0069_ };
  assign _1966_[9] = _0191_ + _0241_;
  assign { _2217_[43:42], _1904_[38:22], _2217_[24:21], _1226_, _2217_[19:0] } = { _2219_[43:31], _2069_[32:23], _1317_, _2069_[21:18], _0545_, _0796_, _0258_, _0232_, _0415_, _1558_, _2219_[9:8], _0284_, _0449_, _1233_, _0021_, _0134_, _0324_, _0165_, _1371_ } + { _1942_[86:58], _0905_, _1170_, _2218_[12:1], _0563_ };
  assign _2222_ = { _1334_, _1020_ } + { _0304_, _1166_ };
  assign { _2224_[17:16], _0916_, _2224_[14:0] } = { _2188_[23:19], _0459_, _2188_[17:6] } + { _2064_[11], _1049_, _1566_, _2064_[8:7], _0161_, _1302_, _0870_, _2191_[9:7], _1914_[46:40] };
  assign { _2228_[67:48], _0541_, _2228_[46:41], _1894_[55:48], _2228_[32:27], _1262_, _2228_[25:0] } = { _2014_[16:10], _1988_[54:51], _0291_, _1988_[49], _1383_, _1988_[47:46], _1697_, _1988_[44], _1153_, _1893_[10:7], _1034_, _1893_[5:4], _1374_, _1787_, _0126_, _1328_, _2229_[37:31], _0867_, _0641_, _1752_, _1721_, _1836_, _2229_[25], _0548_, _2015_[20:2], _1369_, _2015_[0], _0799_, _0004_, _1760_ } + { _2198_[35:6], _1443_, _1626_, _0379_, _0019_, _0749_, _0241_, _0140_, _0808_, _1723_, _1245_, _0572_, _2222_, _0254_, _0753_, _1863_, _0166_, _0132_, _1009_, _0483_, _0032_, _0242_, _0166_, _0458_, _1257_, _0748_, _1634_, _1832_, _1760_, _2207_, _0472_, _1619_, _0429_, _0173_ };
  assign { _2230_[12:9], _0078_, _2230_[7:0] } = { _0687_, _1076_, _0560_, _0846_, _0153_, _0600_, _1636_, _0643_, _0843_, _0363_, _0354_, _0531_, _0489_ } + { _2197_[91:90], _0877_, _2197_[88:82], _0599_, _0699_, _0241_ };
  assign _1904_[9:2] = { _0774_, _1037_, _1567_, _0567_, _0975_, _1463_, _0680_, _0289_ } + { _1105_, _0453_, _0071_, _0235_, _0827_, _0575_, _1457_, _0122_ };
  assign { _2199_[27:21], _0996_, _2199_[19:16], _2010_[3:1], _0240_ } = { _2168_[6:1], _0189_, _0993_, _0403_, _0134_, _0893_, _0097_, _0334_, _0661_, _0408_, _0328_ } + { _1972_[22], _1687_, _1972_[20:11], _2112_[42:41], _0206_, _0531_ };
  assign { _2233_[52:1], _0965_ } = { _2161_[11:0], _1878_, _0433_, _0848_, _1299_, _1901_[57:39], _1021_, _2022_[8:6], _1160_, _2022_[4:3], _1069_, _2022_[1:0], _1251_, _0805_, _0296_, _0250_, _0154_, _1595_, _1192_, _0069_ } + { _0324_, _2158_[50:48], _1300_, _2158_[46:40], _1563_, _2158_[38:34], _1489_, _2158_[32:0], _1388_ };
  assign { _1988_[41:38], _0130_, _1988_[36], _0725_, _1988_[34:27], _1406_, _1175_, _1988_[24], _0921_, _1988_[22], _1819_, _1988_[20:19] } = { _2041_[31], _1755_, _2041_[29:27], _0189_, _0082_, _0228_, _0082_, _0529_, _1964_[52], _1795_, _1964_[50:48], _1016_, _1964_[46:45], _0492_, _1964_[43], _1706_, _0071_, _0226_ } + { _0514_, _2031_[21:19], _1887_[16], _2031_[17], _1101_, _1814_, _2031_[14:3], _1509_, _0103_, _0189_ };
  assign { _2235_[66:46], _0516_, _1958_[13:4], _2235_[34:22], _0006_, _2235_[20:0] } = { _2118_[90:30], _0485_, _0150_, _0779_, _0793_, _0549_, _0005_ } + { _2153_[25:24], _1508_, _2153_[22:0], _1005_, _2236_[39:32], _1700_, _2236_[30:25], _1224_, _0664_, _2236_[22:19], _2215_[7:2], _1559_, _2213_[23:18], _2236_[5:4], _2208_[3:1], _1281_ };
  assign { _2238_[122:87], _1522_, _2238_[85:81], _2212_, _2238_[73:72], _0378_, _2238_[70:57], _1673_, _2016_[21:6], _2238_[39:31], _1943_[111], _1768_, _1943_[109:89], _1007_, _2238_[6:5], _1771_, _2238_[3:0] } = { _1989_[30:5], _1792_, _1989_[3:2], _1992_[8], _2168_[56:16], _0609_, _0241_, _0071_, _1900_[72:70], _0389_, _1900_[68:66], _0833_, _1305_, _1900_[63], _1136_, _0752_, _0096_, _0071_, _0193_, _1136_, _1046_, _0359_, _0109_, _1900_[72:70], _0389_, _1900_[68:66], _0833_, _1305_, _1900_[63], _2199_[27:21], _0996_, _2199_[19:16], _2010_[3:1], _0240_, _0197_, _0232_, _0893_, _0194_ } + { _1951_[154:151], _1276_, _1951_[149:144], _1042_, _1951_[142:139], _0124_, _0929_, _1951_[136], _1530_, _0588_, _1890_[11], _0350_, _0716_, _1890_[8:6], _0294_, _0205_, _2000_[123:108], _1361_, _2000_[106:100], _1506_, _2000_[98], _0113_, _2000_[96:92], _0313_, _2000_[90:86], _0737_, _2000_[84:80], _0354_, _0226_, _0071_, _0463_, _0134_, _0043_, _2121_[43:39], _0864_, _1346_, _2121_[36:35], _1600_, _2121_[33:28], _0653_, _2121_[26:22], _2031_[66], _0328_, _2031_[64], _0007_, _1699_, _2031_[61:55], _1806_, _2031_[53], _0206_, _2031_[51], _1800_, _2031_[49:47], _2121_[1:0] };
  reg [12:0] _3618_;
  always_ff @(posedge _0356_, posedge _1225_)
    if (_1225_) _3618_ <= 13'h128f;
    else _3618_ <= { _0120_, _1568_, _1976_[10:9], _0604_, _1976_[7], _0945_, _1976_[5], _0602_, _1976_[3], _0383_, _0134_, _1170_ };
  assign { _0920_, _2004_[10:6], _1387_, _2018_[58:56], _0397_, _1640_, _2018_[53] } = _3618_;
  reg [1:0] _3619_;
  always_ff @(posedge _0254_, negedge _0708_)
    if (!_0708_) _3619_ <= 2'h2;
    else _3619_ <= { _0306_, _1733_ };
  assign _1957_[1:0] = _3619_;
  reg [8:0] _3620_;
  always_ff @(negedge _0926_, negedge _0354_)
    if (!_0354_) _3620_ <= 9'h1a9;
    else _3620_ <= { _0752_, _0159_, _0118_, _1077_, _0248_, _1684_, _2028_[3], _1326_, _2028_[1] };
  assign { _0986_, _1908_[14:13], _1564_, _1908_[11:10], _0535_, _1908_[8:7] } = _3620_;
  reg [12:0] _3621_;
  always_ff @(negedge _0904_, negedge _0609_)
    if (!_0609_) _3621_ <= 13'h06e0;
    else _3621_ <= { _2243_[12:9], _0768_, _0276_, _0116_, _0127_, _1046_, _0626_, _0227_, _1229_, _1518_ };
  assign _1967_[35:23] = _3621_;
  reg [21:0] _3622_;
  always_ff @(negedge _0106_, negedge _0069_)
    if (!_0069_) _3622_ <= 22'h25ff3a;
    else _3622_ <= { _1979_[41:36], _0084_, _0383_, _0920_, _2004_[10:6], _1387_, _2018_[58:56], _0397_, _1640_, _2018_[53], _0521_ };
  assign { _2242_[21], _1316_, _2242_[19:18], _0616_, _2242_[16], _1378_, _2242_[14:1], _1778_ } = _3622_;
  reg [3:0] _3623_;
  always_ff @(negedge _0019_, negedge _2000_[28])
    if (!_2000_[28]) _3623_ <= 4'h9;
    else _3623_ <= { _0359_, _0565_, _0915_, _0197_ };
  assign { _1810_, _0123_, _1932_[6], _0595_ } = _3623_;
  reg [82:0] _3624_;
  always_ff @(negedge _2105_[42], negedge _0356_)
    if (!_0356_) _3624_ <= 83'h000000000000000000000;
    else _3624_ <= { _0049_, _0752_, _1070_, _2245_[79], _1313_, _0624_, _2141_[22:19], _2245_[72:70], _1984_[46:39], _1714_, _1984_[37:36], _0251_, _1984_[34:15], _2245_[37:34], _1922_, _2245_[30:28], _2091_[14:13], _0644_, _2091_[11], _2014_[17:10], _1988_[54:51], _0291_, _1988_[49], _1383_, _1988_[47:46], _1697_, _1988_[44:43], _0228_, _0191_, _0325_, _0453_ };
  assign { _2244_[82:81], _0970_, _2244_[79:67], _1319_, _2244_[65:56], _2059_[95:89], _0992_, _2059_[87:76], _0547_, _2059_[74:71], _1282_, _2059_[69:67], _1608_, _2059_[65:55], _0822_, _2059_[53:44], _2244_[3:0] } = _3624_;
  reg [1:0] _3625_;
  always_ff @(posedge _2037_[75], negedge _1650_)
    if (!_1650_) _3625_ <= 2'h1;
    else _3625_ <= { _0571_, _1598_ };
  assign { _0086_, _2246_[0] } = _3625_;
  reg [41:0] _3626_;
  always_ff @(posedge _1589_, negedge _0118_)
    if (!_0118_) _3626_ <= 42'h3ffa5bcd1a9;
    else _3626_ <= { _1951_[168:159], _1255_, _1951_[157:151], _1276_, _1951_[149:144], _1042_, _1951_[142:139], _0124_, _0929_, _1951_[136:134], _1493_, _2020_[10:9], _0293_, _2020_[7:5] };
  assign { _2142_[45:43], _1830_, _0093_, _2142_[40:28], _1775_, _2142_[26:18], _2032_[66:54], _2142_[4] } = _3626_;
  reg [40:0] _3627_;
  always_ff @(posedge _1376_, negedge _0642_)
    if (!_0642_) _3627_ <= 41'h1ff9dc60d83;
    else _3627_ <= { _1332_, _2170_[24:12], _0250_, _0154_, _0197_, _2242_[21], _1316_, _2242_[19:18], _0616_, _2242_[16], _1378_, _2242_[14:1], _1778_, _0149_, _0044_ };
  assign { _2059_[42:32], _1474_, _2059_[30:23], _1330_, _2059_[21:18], _1382_, _2059_[16:6], _1249_, _2059_[4:2] } = _3627_;
  reg [54:0] _3628_;
  always_ff @(negedge _1655_, posedge _0226_)
    if (_0226_) _3628_ <= 55'h00000036e2b969;
    else _3628_ <= { _2059_[30], _0134_, _0354_, _1203_, _0109_, _1046_, _0221_, _1362_, _1786_, _0402_, _1397_, _1569_, _1970_[5], _0152_, _0014_, _0200_, _0359_, _0071_, _0642_, _0152_, _1009_, _0149_, _0434_, _1589_, _1206_, _0111_, _0014_, _0919_, _0359_, _0464_, _1976_[19:16], _1335_, _1976_[14], _0172_, _0120_, _1568_, _1976_[10:9], _0604_, _1976_[7], _0945_, _1976_[5], _0602_, _1976_[3:0], _0591_, _0356_, _0993_, _0403_, _0277_ };
  assign { _2254_[54:53], _0878_, _2254_[51], _2054_[40:39], _2039_[13:11], _1417_, _2054_[34:31], _1683_, _2054_[29:19], _1538_, _2054_[17:16], _1029_, _2054_[14:9], _2254_[18], _1717_, _2254_[16:14], _1404_, _2254_[12], _1798_, _2254_[10:2], _0167_, _2254_[0] } = _3628_;
  reg [34:0] _3629_;
  always_ff @(posedge _1733_, negedge _1660_)
    if (!_1660_) _3629_ <= 35'h7980ed188;
    else _3629_ <= { _2146_[19:8], _0821_, _0637_, _1399_, _0216_, _1884_, _0727_, _2008_[14:3], _1531_, _1068_, _2008_[0], _1873_, _0469_ };
  assign { _2255_[34:32], out_data[1503:1472] } = _3629_;
  reg [22:0] _3630_;
  always_ff @(negedge _0670_, negedge _1103_)
    if (!_1103_) _3630_ <= 23'h339b31;
    else _3630_ <= { _0678_, _0116_, _0902_, _1772_, _1900_[62:59], _0498_, _1900_[57:54], _0066_, _1900_[52:50], _0542_, _0887_, _0466_, _0489_, _0963_, _0808_ };
  assign out_data[1174:1152] = _3630_;
  reg [22:0] _3631_;
  always_ff @(posedge _2140_[5], negedge _1734_)
    if (!_1734_) _3631_ <= 23'h034824;
    else _3631_ <= { _1953_[24:11], _0761_, _0360_, _0141_, _0259_, _0449_, _1234_, _0931_, _0555_, _0462_ };
  assign out_data[1014:992] = _3631_;
  reg [6:0] _3632_;
  always_ff @(posedge _1436_, negedge _0016_)
    if (!_0016_) _3632_ <= 7'h12;
    else _3632_ <= { _1151_, _1237_, _0702_, _1858_, _0570_, _0687_, _1473_ };
  assign out_data[358:352] = _3632_;
  reg [65:0] _3633_;
  always_ff @(posedge _1170_, negedge _0018_)
    if (!_0018_) _3633_ <= 66'h00000000000000000;
    else _3633_ <= { _1441_, _2095_[117:108], _1972_[25:22], _1687_, _1972_[20:19], _0018_, _0232_, _0661_, _1994_[9:6], _0840_, _1994_[4:3], _0597_, _2048_[51:50], _1423_, _2048_[48:47], _2005_[10:8], _1327_, _2005_[6:4], _2048_[39:38], _1150_, _2048_[36], _1010_, _2048_[34:17], _0226_, _0277_ };
  assign { _2256_[65:49], _1969_[51:36], _0677_, _1969_[34:29], _0985_, _1969_[27:8], _2256_[4:0] } = _3633_;
  reg [36:0] _3634_;
  always_ff @(posedge _1018_, negedge _0820_)
    if (!_0820_) _3634_ <= 37'h1fefe4d83f;
    else _3634_ <= { _1169_, _1176_, _1557_, _1956_[30:24], _1618_, _1956_[22], _2140_[13:0], _1962_[11:5], _1261_, _1962_[3:1] };
  assign { _2257_[36], out_data[63:32], _2257_[3:0] } = _3634_;
  reg [59:0] _3635_;
  always_ff @(negedge _0177_, negedge _0922_)
    if (!_0922_) _3635_ <= 60'hfffffffda06d234;
    else _3635_ <= { _2170_[32:31], _1008_, _2170_[29:26], _1332_, _2170_[24:19], _1374_, _1266_, _2000_[123:108], _1361_, _2000_[106:100], _1506_, _2000_[98], _0113_, _2000_[96:92], _0313_, _2000_[90:86], _0737_, _2000_[84:80] };
  assign { _2001_[139:138], _0211_, _2001_[136:113], _2234_[21:6], _2132_[1], _0791_, _2258_[14:0] } = _3635_;
  reg [47:0] _3636_;
  always_ff @(posedge _0059_, posedge _0082_)
    if (_0082_) _3636_ <= 48'h000058536e2f;
    else _3636_ <= { _2121_[41:39], _0864_, _1346_, _2121_[36:35], _1600_, _2121_[33:28], _0653_, _2121_[26:22], _2031_[66], _0328_, _2031_[64], _0007_, _1699_, _2031_[61:55], _1806_, _2031_[53], _0206_, _2031_[51], _1800_, _2031_[49:47], _0408_, _0311_, _0490_, _0044_, _0270_, _0304_, _0636_, _0661_ };
  assign { _1976_[70:58], _1797_, _1976_[56:34], _0100_, _1976_[32:26], _1341_, _1976_[24:23] } = _3636_;
  reg [24:0] _3637_;
  always_ff @(negedge _1381_, posedge _1009_)
    if (_1009_) _3637_ <= 25'h0fa2f32;
    else _3637_ <= { _1971_[24:19], _0922_, _1971_[17:13], _1525_, _1971_[11:1], _0924_ };
  assign { _2001_[95:86], _0998_, _2001_[84:73], _1765_, _2001_[71] } = _3637_;
  reg [7:0] _3638_;
  always_ff @(negedge _1970_[5], negedge _1346_)
    if (!_1346_) _3638_ <= 8'h0d;
    else _3638_ <= { _1972_[11], _2112_[42:40], _0191_, _0097_, _0150_, _0071_ };
  assign { _1866_, _2225_[10], _0962_, _2225_[8:4] } = _3638_;
  reg [25:0] _3639_;
  always_ff @(negedge _0152_, posedge _0359_)
    if (_0359_) _3639_ <= 26'h29acd34;
    else _3639_ <= { _1969_[30:29], _0985_, _1969_[27:15], _0149_, _0482_, _1761_, _1590_, _1929_[4:3], _0103_, _0453_, _0524_, _0591_ };
  assign { _1966_[39:34], _0990_, _1966_[32:27], _0988_, _1879_, _1966_[24:19], _0528_, _1966_[17:14] } = _3639_;
  reg [37:0] _3640_;
  always_ff @(posedge _0919_, posedge _0227_)
    if (_0227_) _3640_ <= 38'h0010e2e9e8;
    else _3640_ <= { _2244_[65:56], _2059_[95:93], _0159_, _0038_, _2242_[21], _1316_, _2242_[19:18], _0616_, _2242_[16], _1378_, _2242_[14:1], _1778_, _0453_ };
  assign { _2108_[80:78], _1791_, _2108_[76], _2053_[40:28], _1667_, _2053_[26:21], _1695_, _2053_[19:15], _1185_, _2053_[13:11], _2108_[45:43] } = _3640_;
  reg [53:0] _3641_;
  always_ff @(posedge _0243_, posedge _0099_)
    if (_0099_) _3641_ <= 54'h3fffffb5342b63;
    else _3641_ <= { _0502_, _0058_, _0197_, _1994_[9:6], _0840_, _1994_[4:3], _0597_, _2048_[51:50], _1423_, _2048_[48:47], _2005_[10:8], _1327_, _2005_[6:4], _2048_[39:38], _1150_, _2048_[36], _1010_, _2048_[34:17], _0102_, _0134_, _1014_, _1952_[141], _1621_, _1577_, _1320_, _1952_[137] };
  assign { _2219_[43:31], _2069_[32:23], _1317_, _2069_[21:13], _2259_[20:19], _2085_[9], _2074_[6], _2049_[83:72], _1121_, _2049_[70:69], _1670_, _2259_[0] } = _3641_;
  reg [3:0] _3642_;
  always_ff @(posedge _0593_, negedge _0108_)
    if (!_0108_) _3642_ <= 4'hf;
    else _3642_ <= { _2238_[100:98], _0044_ };
  assign { _1951_[33], _1412_, _1951_[31], _1496_ } = _3642_;
  reg [53:0] _3643_;
  always_ff @(posedge _0893_, negedge _2040_[18])
    if (!_2040_[18]) _3643_ <= 54'h00000000c2ce14;
    else _3643_ <= { _2242_[7], _0299_, _0275_, _0563_, _1983_[46:26], _1928_[24:18], _0244_, _1928_[16:12], _0441_, _1928_[10:9], _1983_[9:0], _0151_, _1000_, _0287_ };
  assign { _2019_[58:57], _1636_, _2019_[55:37], _0070_, _1920_[31:22], _0056_, _1920_[20:19], _1816_, _1920_[17:16], _1168_, _1920_[14:2], _2019_[5] } = _3643_;
  reg [15:0] _3644_;
  always_ff @(posedge _1971_[15], negedge _2025_[32])
    if (!_2025_[32]) _3644_ <= 16'h07f3;
    else _3644_ <= { _0364_, _1888_[13], _0036_, _0706_, _1888_[10:5], _0673_, _1964_[55], _0983_, _0354_, _0134_, _0254_ };
  assign { _2139_[66:60], _1705_, _2139_[58:55], _1743_, _0943_, _2139_[52:51] } = _3644_;
  reg [8:0] _3645_;
  always_ff @(posedge _0238_, negedge _0082_)
    if (!_0082_) _3645_ <= 9'h013;
    else _3645_ <= { _2053_[32:28], _1667_, _2053_[26:24] };
  assign { _1337_, _2054_[7:2], _1633_, _0156_ } = _3645_;
  reg [21:0] _3646_;
  always_ff @(negedge _0210_, posedge _1951_[31])
    if (_1951_[31]) _3646_ <= 22'h23ba6e;
    else _3646_ <= { _2244_[71:70], _0748_, _0152_, _0915_, _1956_[18:15], _0506_, _1956_[13:12], _0591_, _0096_, _0600_, _0082_, _0617_, _0566_, _0238_, _0189_, _1283_, _1113_ };
  assign { _1967_[21:15], _1668_, _1967_[13:10], _1321_, _0473_, _1967_[7:0] } = _3646_;
  reg [11:0] _3647_;
  always_ff @(negedge _0241_, negedge _0356_)
    if (!_0356_) _3647_ <= 12'h653;
    else _3647_ <= { _2095_[114:112], _0200_, _0356_, _0043_, _0250_, _0154_, _0359_, _0226_, _0025_, _0152_ };
  assign { _1153_, _1893_[10:7], _1034_, _1893_[5:4], _1374_, _1787_, _0126_, _1328_ } = _3647_;
  reg [25:0] _3648_;
  always_ff @(posedge _1323_, negedge _0049_)
    if (!_0049_) _3648_ <= 26'h1df14df;
    else _3648_ <= { _2238_[88:87], _1522_, _2238_[85:81], _2212_, _2238_[73:72], _0378_, _2238_[70:67], _0638_, _0984_, _0316_, _0477_ };
  assign { _2064_[37], _1350_, _2064_[35:34], _2024_[13:12], _1825_, _2024_[10:2], _2064_[21:14], _1676_, _2064_[12] } = _3648_;
  reg [36:0] _3649_;
  always_ff @(posedge _1939_[10], posedge _1564_)
    if (_1564_) _3649_ <= 37'h1fc8d0d924;
    else _3649_ <= { _2000_[15:14], _0925_, _1939_[12:11], _0165_, _0071_, _0134_, _0221_, _0356_, _2000_[20:19], _0564_, _2000_[17:14], _0925_, _1939_[12:8], _0501_, _1939_[6], _1306_, _2000_[4:3], _1632_, _1373_, _2000_[0], _0146_, _0113_, _1632_, _0572_, _0238_, _0044_ };
  assign { _1943_[37:25], _1498_, _1943_[23:5], _0647_, _1943_[3:1] } = _3649_;
  reg [34:0] _3650_;
  always_ff @(posedge _2203_[2], negedge _0154_)
    if (!_0154_) _3650_ <= 35'h7eba1c50f;
    else _3650_ <= { _2053_[25:21], _1695_, _2053_[19:15], _1185_, _2053_[13:11], _2108_[45:43], _0208_, _0354_, _1964_[67], _0364_, _1888_[13], _0036_, _0706_, _1888_[10:5], _0673_, _1964_[55], _1679_, _1170_ };
  assign { _2119_[37:30], _1450_, _1638_, _2119_[27:26], _1502_, _2119_[24:20], _0828_, _2051_[9], _2119_[17], _1106_, _2119_[15:14], _1171_, _2119_[12:3] } = _3650_;
  reg [66:0] _3651_;
  always_ff @(negedge _2112_[35], posedge in_data[767])
    if (in_data[767]) _3651_ <= 67'h00000000035c378db;
    else _3651_ <= { in_data[609:547], _0127_, _0043_, _0096_, _0132_ };
  assign { _2169_[101], _2105_[43:38], _2035_[23:19], _1455_, _1507_, _2035_[16], _1674_, _2035_[14:2], _2082_[30:27], _0628_, _2082_[25:24], _1223_, _2082_[22:19], _1355_, _2082_[17:15], _2169_[56:55], _0451_, _2169_[53:45], _1793_, _2169_[43:40], _1324_, _2169_[38:35] } = _3651_;
  reg [42:0] _3652_;
  always_ff @(posedge _2040_[19], negedge _0379_)
    if (!_0379_) _3652_ <= 43'h0003a4f2fa2;
    else _3652_ <= { _2000_[20:19], _0564_, _2000_[17:14], _0925_, _1939_[12:8], _0501_, _1939_[6], _1956_[18:15], _0506_, _1956_[13:12], _0174_, _1310_, _1393_, _0983_, _0463_, _0194_, _0206_, _1493_, _2020_[10:9], _0293_, _2020_[7:5], _1632_, _0189_, _0144_, _0317_, _0502_, _0095_, _0191_ };
  assign { _2260_[42:23], _2056_[3:1], _2260_[19:13], _0806_, _2260_[11:0] } = _3652_;
  reg [109:0] _3653_;
  always_ff @(posedge _0058_, negedge _1302_)
    if (!_1302_) _3653_ <= 110'h0000000000000000000000000000;
    else _3653_ <= { _0597_, _2048_[51:50], _1423_, _2048_[48:47], _2005_[10:8], _1327_, _2005_[6:4], _2048_[39:38], _1150_, _2048_[36], _1010_, _2048_[34:28], _0477_, _0651_, _0163_, _1203_, _0522_, _1206_, _1113_, _0408_, _0811_, _1956_[18:15], _0506_, _1956_[13:12], _0591_, _0795_, _0275_, _0887_, _0110_, _0334_, _0926_, _0674_, _0610_, _2067_[2:1], _0775_, _2262_[56:54], _1690_, _2262_[52], _2025_[43:40], _1785_, _2025_[38:34], _1510_, _2025_[32:27], _0896_, _2025_[25], _1556_, _0114_, _0319_, _2041_[32:31], _1755_, _2041_[29:24], _0233_, _0499_, _2114_[25:23], _0071_, _1964_[67], _0364_, _1888_[13], _0036_, _0706_, _1888_[10:5], _0673_, _1964_[55], _1679_, _1311_ };
  assign { _2261_[109:104], _1104_, _2261_[102:68], _2026_[43:34], _0842_, _2026_[32:11], _1097_, _2026_[9:7], _2261_[30:26], _1045_, _2261_[24:0] } = _3653_;
  reg [9:0] _3654_;
  always_ff @(negedge _0524_, posedge _0185_)
    if (_0185_) _3654_ <= 10'h32f;
    else _3654_ <= { _1991_[49:47], _1193_, _1553_, _1991_[44:43], _2031_[33:31] };
  assign { _2139_[49], _1748_, _2139_[47:45], _1837_, _2139_[43], _1256_, _2139_[41:40] } = _3654_;
  reg [59:0] _3655_;
  always_ff @(posedge _1203_, negedge _0391_)
    if (!_0391_) _3655_ <= 60'hfffffffa0b72fed;
    else _3655_ <= { _2019_[50:38], _0049_, _0203_, _0586_, _1998_[40:30], _1325_, _1998_[28:0], _0317_, _0098_, _0272_ };
  assign { _2101_[165:163], _2045_[8:5], _2012_[43:28], _1625_, _2012_[26:22], _1678_, _1222_, _2012_[19:2], _1613_, _2101_[115:111], _2263_[4:0] } = _3655_;
  reg [1:0] _3656_;
  always_ff @(negedge _0013_, negedge _0117_)
    if (!_0117_) _3656_ <= 2'h0;
    else _3656_ <= { _0019_, _1393_ };
  assign { _1396_, _1131_ } = _3656_;
  reg [90:0] _3657_;
  always_ff @(posedge _1974_[0], posedge _0617_)
    if (_0617_) _3657_ <= 91'h00000000000000000000000;
    else _3657_ <= { _1795_, _1964_[50:48], _1016_, _1964_[46], _0278_, _0334_, _0140_, _0134_, _0335_, _1786_, _0402_, _1397_, _1569_, _1970_[5], _1493_, _2020_[10:9], _0293_, _2020_[7:5], _1136_, _0221_, _0146_, _0210_, _0748_, _1235_, _1247_, _0549_, _0096_, _0251_, _1337_, _2054_[7:2], _1633_, _0156_, _0145_, _0572_, _0189_, _0042_, _0856_, _2121_[43:39], _0864_, _1346_, _2121_[36:35], _1600_, _2121_[33:28], _0653_, _2121_[26:22], _2031_[66], _0328_, _2031_[64], _0007_, _1699_, _2031_[61:55], _1806_, _2031_[53], _0206_, _2031_[51], _1800_, _2031_[49:47], _2121_[1:0] };
  assign { _1503_, _2111_[50:35], _2264_[73:59], _0968_, _2264_[57:52], _1802_, _2264_[50:17], _2043_[12:2], _2264_[5:0] } = _3657_;
  reg [8:0] _3658_;
  always_ff @(posedge _2026_[36], posedge _0254_)
    if (_0254_) _3658_ <= 9'h110;
    else _3658_ <= { _2059_[10:9], _0059_, _0633_, _0162_, _1959_[7], _1202_, _0016_, _0238_ };
  assign { _2022_[8:6], _1160_, _2022_[4:3], _1069_, _2022_[1:0] } = _3658_;
  reg [1:0] _3659_;
  always_ff @(posedge _0025_, negedge _0025_)
    if (!_0025_) _3659_ <= 2'h1;
    else _3659_ <= { _0200_, _0025_ };
  assign { _0250_, _0154_ } = _3659_;
  reg [17:0] _3660_;
  always_ff @(negedge _0134_, posedge _2169_[38])
    if (_2169_[38]) _3660_ <= 18'h36b4f;
    else _3660_ <= { _2006_[6], _0404_, _2006_[4:3], _1931_[3], _1308_, _0513_, _1254_, _0468_, _2006_[6], _0404_, _2006_[4:3], _1931_[3], _1308_, _0513_, _0359_, _0033_ };
  assign { _2040_[20:11], _0618_, _1485_, _2040_[8], _1488_, _2040_[6:3] } = _3660_;
  reg [61:0] _3661_;
  always_ff @(posedge _0626_, posedge _1381_)
    if (_1381_) _3661_ <= 62'h000000002f1522bc;
    else _3661_ <= { _2216_[87:86], _0734_, _0306_, _0211_, _0024_, _0589_, _0469_, _0128_, out_data[416], _0096_, _0204_, _0134_, _2119_[37:30], _1450_, _1638_, _2119_[27:26], _1502_, _2119_[24:20], _0828_, _2051_[9], _2119_[17], _1106_, _2119_[15:14], _1171_, _2119_[12:3], _0092_, _0254_, _1993_[9:6], _1041_, _1993_[4:0], _0598_, _0318_ };
  assign { _2265_[61:48], _1333_, _2265_[46:38], _2241_[39], _1936_[79:55], _2241_[13:4], _2265_[1:0] } = _3661_;
  reg [1:0] _3662_;
  always_ff @(negedge _0620_, posedge _0989_)
    if (_0989_) _3662_ <= 2'h3;
    else _3662_ <= _2006_[4:3];
  assign { _1836_, _2229_[25] } = _3662_;
  reg [8:0] _3663_;
  always_ff @(posedge _0361_, posedge _0320_)
    if (_0320_) _3663_ <= 9'h003;
    else _3663_ <= { in_data[1882:1879], _0907_, _0854_, _0149_, _0071_, _0025_ };
  assign { _1846_, _1248_, _2231_[159], _0045_, _2231_[157:156], _1751_, _1536_, _2231_[153] } = _3663_;
  reg [104:0] _3664_;
  always_ff @(posedge _0113_, posedge _0146_)
    if (_0146_) _3664_ <= 105'h000000000000000000000000000;
    else _3664_ <= { in_data[1797:1746], _0733_, _0140_, _1014_, _1952_[141], _1621_, _1577_, _1320_, _1952_[137], _0270_, _0565_, _0251_, _2164_[29:24], _0601_, _2164_[22:20], _1997_, _2164_[16:12], _2154_[39:35], _1080_, _2154_[33:32], _1338_, _2164_[2:0], _1981_[11:9], _0299_, _0223_, _1981_[6:2], _1794_, _0140_ };
  assign { _2266_[104:96], _2183_[102:50], _1349_, _2183_[48:29], _2079_[21:4], _2266_[3:0] } = _3664_;
  reg [44:0] _3665_;
  always_ff @(posedge _0469_, negedge _0016_)
    if (!_0016_) _3665_ <= 45'h0000741e2679;
    else _3665_ <= { _1983_[43:26], _1928_[24:18], _0244_, _1928_[16:12], _0068_, _0116_, _0311_, _0052_, _0197_, _0103_, _0151_, _0984_, _0127_, _1211_, _0134_, _0141_, _1449_, _1552_ };
  assign { _2038_[44:43], _0630_, _0407_, _2038_[40:25], _1060_, _2038_[23:11], _2034_[23:15], _2038_[1:0] } = _3665_;
  always_ff @(negedge _0165_, negedge _0748_)
    if (!_0748_) _0380_ <= 1'h0;
    else _0380_ <= _1787_;
  reg [10:0] _3667_;
  always_ff @(posedge _0065_, posedge _0359_)
    if (_0359_) _3667_ <= 11'h7c5;
    else _3667_ <= { _1990_[8:1], _0018_, _0593_, _0726_ };
  assign { _2267_[10:7], _1214_, _2267_[5:0] } = _3667_;
  reg [98:0] _3668_;
  always_ff @(posedge _0226_, negedge _0549_)
    if (!_0549_) _3668_ <= 99'h0000000000000000000000000;
    else _3668_ <= { _1976_[66:58], _1797_, _1976_[56:43], _0237_, _0189_, _1072_, _0453_, _0325_, _0254_, _1134_, _0609_, _0227_, _2000_[59:50], _1570_, _2000_[48:46], _1314_, _1419_, _0391_, _2000_[42:35], _1747_, _2000_[33:31], _1307_, _2000_[29:27], _1318_, _0228_, _2267_[10:7], _1214_, _2267_[5:0], _0361_, _0334_, _1206_, _0748_, _0254_, _0043_, _0726_, _0092_, _0105_, _0452_, _0469_, _0572_, _0642_, _0524_, _0096_, _0116_, _0590_, _0603_, _0598_, _0254_ };
  assign { _2268_[98:78], _1961_[34:1], _2268_[43:38], _2038_[80:48], _1039_, _2038_[46], _2268_[2:0] } = _3668_;
  reg [1:0] _3669_;
  always_ff @(posedge _0586_, negedge _0134_)
    if (!_0134_) _3669_ <= 2'h2;
    else _3669_ <= { _0101_, _0200_ };
  assign { _0081_, _1340_ } = _3669_;
  reg [32:0] _3670_;
  always_ff @(negedge _1211_, negedge _1982_[13])
    if (!_1982_[13]) _3670_ <= 33'h01f530467;
    else _3670_ <= { _2025_[40], _1785_, _2025_[38:34], _1510_, _2025_[32:27], _0896_, _2025_[25], _1556_, _0114_, _0319_, _2041_[32:31], _1755_, _2041_[29:24], _0233_, _0499_, _2114_[25:23] };
  assign { _2245_[36:34], _1922_, _2245_[30:28], _2091_[14:13], _0644_, _2091_[11], _2014_[17:10], _1988_[54:51], _0291_, _1988_[49], _1383_, _1988_[47:46], _1697_, _1988_[44:43] } = _3670_;
  reg [2:0] _3671_;
  always_ff @(negedge _0259_, negedge _0272_)
    if (!_0272_) _3671_ <= 3'h1;
    else _3671_ <= { _0019_, _0490_, _0995_ };
  assign { _1893_[50:49], _0771_ } = _3671_;
  always_ff @(posedge _0739_, posedge _2059_[7])
    if (_2059_[7]) _1360_ <= 1'h1;
    else _1360_ <= _0733_;
  reg [3:0] _3673_;
  always_ff @(negedge _2012_[23], negedge _0254_)
    if (!_0254_) _3673_ <= 4'ha;
    else _3673_ <= { _1995_[6], _1242_, _1086_, _0678_ };
  assign { _1935_[18:17], _0558_, _1935_[15] } = _3673_;
  reg [8:0] _3674_;
  always_ff @(posedge _0117_, posedge _0748_)
    if (_0748_) _3674_ <= 9'h0df;
    else _3674_ <= _1984_[24:16];
  assign { _2139_[35:32], _1354_, _1054_, _2139_[29:27] } = _3674_;
  reg [6:0] _3675_;
  always_ff @(negedge _0354_, negedge _1997_[0])
    if (!_1997_[0]) _3675_ <= 7'h71;
    else _3675_ <= { _2139_[49], _1748_, _2139_[47], _0259_, _0380_, _0116_, _0016_ };
  assign { _2046_[6], _1756_, _2046_[4], _1094_, _2046_[2:0] } = _3675_;
  reg [4:0] _3676_;
  always_ff @(negedge _2022_[1], posedge _1909_[12])
    if (_1909_[12]) _3676_ <= 5'h1c;
    else _3676_ <= { _1976_[16], _1335_, _1976_[14], _0172_, _0120_ };
  assign { _2220_[17:15], _1032_, _2220_[13] } = _3676_;
  reg [11:0] _3677_;
  always_ff @(posedge _0455_, posedge _1004_)
    if (_1004_) _3677_ <= 12'h28d;
    else _3677_ <= { _2001_[104:103], _1351_, _2001_[101], _0936_, _0163_, _0994_, _1391_, _0143_, _0299_, _0092_, _0984_ };
  assign { _1955_[25:20], _0072_, _1955_[18], _1853_, _1955_[16], _1487_, _1955_[14] } = _3677_;
  reg [12:0] _3678_;
  always_ff @(negedge _0102_, posedge _2267_[10])
    if (_2267_[10]) _3678_ <= 13'h1606;
    else _3678_ <= { _1980_[13:10], _0299_, _0258_, _0648_, _0272_, _2220_[17:15], _1032_, _2220_[13] };
  assign { _2269_[12], _0892_, _2269_[10:8], _1050_, _0329_, _1813_, _2269_[4:0] } = _3678_;
  reg [76:0] _3679_;
  always_ff @(negedge _0108_, posedge _2059_[60])
    if (_2059_[60]) _3679_ <= 77'h00000000000000000000;
    else _3679_ <= { _1912_[29:24], _0781_, _1994_[9:6], _0840_, _1994_[4:3], _0597_, _2048_[51:50], _1423_, _2048_[48:47], _2005_[10:8], _1327_, _2005_[6:4], _2048_[39:38], _1150_, _2048_[36], _1010_, _2048_[34:17], _0152_, _0633_, _0162_, _1959_[7], _1202_, _0857_, _0420_, _0062_, _0793_, _1464_, _2022_[8:6], _1160_, _2022_[4:3], _1069_, _2022_[1:0], _1956_[18:15], _0506_, _1956_[13:12], _0893_ };
  assign { _2270_[76:67], _0667_, _2094_[130:103], _1291_, _2094_[101:94], _1263_, _2094_[92:69], _2270_[3:0] } = _3679_;
  reg [48:0] _3680_;
  always_ff @(negedge _0357_, negedge _0097_)
    if (!_0097_) _3680_ <= 49'h000000def156e;
    else _3680_ <= { _1034_, _1893_[5], _1000_, _0096_, _2032_[31:26], _1826_, _2032_[24:13], _0606_, _2032_[11:10], _1754_, _2032_[8:1], _1551_, _1846_, _1248_, _2231_[159], _0045_, _2231_[157:156], _1751_, _1536_, _2231_[153], _0795_, _0755_, _0228_, _0194_ };
  assign { _2271_[48:38], _1694_, _2271_[36:0] } = _3680_;
  reg [23:0] _3681_;
  always_ff @(negedge _1493_, negedge _0116_)
    if (!_0116_) _3681_ <= 24'h9a3e7f;
    else _3681_ <= { _1982_[21:16], _1534_, _1982_[14:6], _1287_, _2002_[6:5], _1551_, _0454_, _0678_, _0589_, _0452_ };
  assign { _2272_[23:15], _2252_, _2272_[13], _2104_[6:3], _2272_[8:0] } = _3681_;
  reg [22:0] _3682_;
  always_ff @(posedge _0076_, negedge _0217_)
    if (!_0217_) _3682_ <= 23'h2683b4;
    else _3682_ <= { _2001_[111], _1323_, _2001_[109], _1309_, _1081_, _2001_[106:103], _1351_, _2001_[101:100], _0987_, _1552_, _1254_, _0468_, _2006_[6], _0404_, _2006_[4:3], _1931_[3], _1308_, _0513_ };
  assign { _1898_[38:23], _1517_, _1898_[21:17], _1593_ } = _3682_;
  reg [69:0] _3683_;
  always_ff @(negedge _2183_[91], negedge _0697_)
    if (!_0697_) _3683_ <= 70'h000000000000000000;
    else _3683_ <= { _2017_[65:61], _1364_, _2017_[59:37], _1410_, _2017_[35:33], _0414_, _2017_[31:14], _1442_, _2017_[12:0], _0272_, _1056_, _0609_, _0118_ };
  assign { _2273_[69:28], _1919_[31:17], _0557_, _1919_[15:7], _1882_, _1919_[5], _2273_[0] } = _3683_;
  reg [20:0] _3684_;
  always_ff @(posedge _0315_, posedge _0053_)
    if (_0053_) _3684_ <= 21'h024fb7;
    else _3684_ <= { _1976_[18:16], _1335_, _1976_[14], _0172_, _0120_, _1568_, _1976_[10:9], _0604_, _1976_[7], _0945_, _1976_[5], _0602_, _1976_[3:0], _0608_, _0278_ };
  assign { _2101_[46:40], _1163_, _2101_[38:34], _1216_, _2101_[32:27], _0658_ } = _3684_;
  reg [33:0] _3685_;
  always_ff @(negedge _0133_, posedge _0134_)
    if (_0134_) _3685_ <= 34'h0079f60e7;
    else _3685_ <= { _2003_[9], _1126_, _1631_, _2003_[6:3], _1372_, _0594_, _0920_, _2004_[10:6], _1387_, _2018_[58:56], _0397_, _1640_, _2018_[53], _0643_, _0192_, _0062_, _0096_, _0652_, _1170_, _1561_, _0631_, _0748_, _0024_, _1485_, _0309_ };
  assign { _2274_[33:32], _2209_[32], _0972_, _2201_[12], _2209_[29:16], _1620_, _2209_[14], _1966_[77:65] } = _3685_;
  reg [2:0] _3686_;
  always_ff @(negedge _0434_, posedge _0317_)
    if (_0317_) _3686_ <= 3'h6;
    else _3686_ <= { _1981_[2], _1794_, _0385_ };
  assign { _1579_, _1573_, _2190_[74] } = _3686_;
  reg [18:0] _3687_;
  always_ff @(negedge _0619_, posedge _0215_)
    if (_0215_) _3687_ <= 19'h2423a;
    else _3687_ <= { _2139_[35:32], _1354_, _1054_, _2139_[29:27], _1006_, _0460_, _0166_, _0264_, _0315_, _1627_, _0631_, _1019_, _1130_, _0354_ };
  assign { _2060_[58:51], _0862_, _2060_[49], _2057_[2:1], _2060_[46], _1719_, _2060_[44:40] } = _3687_;
  reg [16:0] _3688_;
  always_ff @(posedge _1751_, negedge _0187_)
    if (!_0187_) _3688_ <= 17'h13a0f;
    else _3688_ <= { _2007_[1], _1441_, _2095_[117:113], _1310_, _0175_, _0283_, _1810_, _0123_, _1932_[6], _0595_, _0111_, _0795_, _0058_ };
  assign { _1468_, _2098_[18:3] } = _3688_;
  reg [2:0] _3689_;
  always_ff @(negedge _1348_, negedge _1339_)
    if (!_1339_) _3689_ <= 3'h4;
    else _3689_ <= { _0401_, _0041_, _1302_ };
  assign _1951_[130:128] = _3689_;
  reg [7:0] _3690_;
  always_ff @(posedge _0594_, posedge _0146_)
    if (_0146_) _3690_ <= 8'hc1;
    else _3690_ <= { _1955_[24:20], _0072_, _1955_[18], _1853_ };
  assign { _1894_[45:41], _0676_, _1894_[39:38] } = _3690_;
  reg [2:0] _3691_;
  always_ff @(negedge _0000_, negedge _1206_)
    if (!_1206_) _3691_ <= 3'h2;
    else _3691_ <= { _1374_, _1787_, _0126_ };
  assign { _1558_, _2219_[9:8] } = _3691_;
  always_ff @(negedge _0109_, negedge _0343_)
    if (!_0343_) _2275_ <= 14'h155c;
    else _2275_ <= { _2069_[27:23], _1317_, _2069_[21:19], _0144_, _0502_, _0041_, _0401_, _0174_ };
  reg [4:0] _3693_;
  always_ff @(posedge _0199_, negedge _1322_)
    if (!_1322_) _3693_ <= 5'h15;
    else _3693_ <= { _0482_, _1761_, _1590_, _1929_[4:3] };
  assign { _2064_[11], _1049_, _1566_, _2064_[8:7] } = _3693_;
  reg [29:0] _3694_;
  always_ff @(negedge _0632_, negedge _0055_)
    if (!_0055_) _3694_ <= 30'h24e5a97c;
    else _3694_ <= { _1981_[11:9], _0299_, _1558_, _2219_[9:8], _0632_, _1639_, _1900_[46:37], _0767_, _1900_[35:29], _0230_, _1833_, _1900_[26] };
  assign { _2111_[33:29], _2087_[31], _2111_[27:21], _1200_, _2111_[19:4] } = _3694_;
  reg [6:0] _3695_;
  always_ff @(negedge _0469_, posedge _0015_)
    if (_0015_) _3695_ <= 7'h12;
    else _3695_ <= { _1007_, _1315_, _0084_, _0420_, _0936_, _1144_, _0463_ };
  assign { _2069_[8], _1458_, _2069_[6:5], _0696_, _1649_, _2069_[2] } = _3695_;
  reg [53:0] _3696_;
  always_ff @(negedge _0235_, posedge _0592_)
    if (_0592_) _3696_ <= 54'h3fffff9b0abc3e;
    else _3696_ <= { _1522_, _2238_[85:81], _2212_, _2238_[73:72], _0378_, _2238_[70:58], _0454_, _0408_, _0343_, _0242_, _0278_, _1809_, _0185_, _0537_, _0481_, _0550_, _0145_, _1981_[11:9], _0299_, _0223_, _1981_[6:2], _1794_, _0521_, _0438_, _0069_ };
  assign { _2223_[55:43], _1896_[35:24], _1594_, _1896_[22:12], _1712_, _1896_[10:9], _2223_[15:2] } = _3696_;
  reg [14:0] _3697_;
  always_ff @(posedge _2069_[28], negedge _0264_)
    if (!_0264_) _3697_ <= 15'h1959;
    else _3697_ <= { _2267_[10:7], _1214_, _2267_[5:2], _0143_, _1966_[4], _0818_, _1966_[2], _0502_, _0748_ };
  assign { _2095_[24], _1661_, _1710_, _2095_[21], _1162_, _1272_, _2095_[18:12], _1585_, _0746_ } = _3697_;
  reg [64:0] _3698_;
  always_ff @(negedge _0590_, posedge _2277_)
    if (_2277_) _3698_ <= 65'h00000000000000000;
    else _3698_ <= { _2030_[54:46], _0705_, _2030_[44:42], _1598_, _2030_[40:16], _1685_, _2030_[14:9], _1468_, _2098_[18:3], _0134_, _0503_ };
  assign { _2276_[64:52], _1637_, _2276_[50:40], _2123_[22:1], _2276_[17:15], _1860_, _2276_[13:0] } = _3698_;
  reg [56:0] _3699_;
  always_ff @(posedge _0032_, posedge _0096_)
    if (_0096_) _3699_ <= 57'h1ffffffcd1c3757;
    else _3699_ <= { _2047_[27:14], _0098_, _0044_, _1998_[40:30], _1325_, _1998_[28:0] };
  assign { _2185_[56:32], _2176_, _1475_, _2185_[22:6], _1703_, _2185_[4:0] } = _3699_;
  reg [56:0] _3700_;
  always_ff @(posedge _0041_, posedge _0566_)
    if (_0566_) _3700_ <= 57'h0000000058b01a1;
    else _3700_ <= { _2029_[40:30], _1012_, _2029_[28:19], _1357_, _2029_[17], _0632_, _1677_, _0409_, _1804_, _1386_, _2002_[27:26], _1381_, _1520_, _1982_[21:16], _1534_, _1982_[14:6], _1287_, _2002_[6:0] };
  assign { _1886_[16], _2278_[55:36], _1738_, _2278_[34:32], out_data[1600], _2278_[30:0] } = _3700_;
  reg [80:0] _3701_;
  always_ff @(negedge _0359_, posedge _0317_)
    if (_0317_) _3701_ <= 81'h000000000000000000000;
    else _3701_ <= { _2082_[28:27], _0628_, _2082_[25:24], _1223_, _2082_[22:19], _1355_, _2082_[17:15], _2169_[56:55], _0451_, _2169_[53:45], _0132_, _0106_, _0189_, _1235_, _0152_, _0068_, _0915_, _0189_, _0084_, _0149_, _2121_[43:39], _0864_, _1346_, _2121_[36:35], _1600_, _2121_[33:28], _0653_, _2121_[26:22], _2031_[66], _0328_, _2031_[64], _0007_, _1699_, _2031_[61:55], _1806_, _2031_[53], _0206_, _2031_[51], _1800_, _2031_[49:47], _2121_[1:0], _0306_ };
  assign { _2170_[84:70], _2070_[32:18], _1201_, _2070_[16:11], _1796_, _2070_[9:5], _0165_, _2070_[3:1], _2170_[37:31], _1008_, _2170_[29:26], _1332_, _2170_[24:9], _0169_, _2170_[7:4] } = _3701_;
  reg [11:0] _3702_;
  always_ff @(negedge _0595_, posedge _2069_[8])
    if (_2069_[8]) _3702_ <= 12'h403;
    else _3702_ <= { _2164_[13:12], _2154_[39:35], _1080_, _1632_, _0209_, _0200_, _1005_ };
  assign _2218_[12:1] = _3702_;
  reg [55:0] _3703_;
  always_ff @(posedge _1331_, negedge _0071_)
    if (!_0071_) _3703_ <= 56'h00000061c073b1;
    else _3703_ <= { _2112_[83:81], _2095_[130:127], _2007_[8:1], _1441_, _2095_[117:108], _1972_[25:22], _1687_, _1972_[20], _0907_, _0702_, _0994_, _0118_, _1015_, _0161_, _2027_[10:9], _0889_, _2027_[7:5], _0260_, _2027_[3:1], _1107_, _0677_, _1027_, _0231_, _0315_, _0690_, _0170_, _1585_ };
  assign { _2279_[55:42], _2083_[28:7], _2279_[19:5], _0556_, _2279_[3:0] } = _3703_;
  reg [5:0] _3704_;
  always_ff @(negedge _0154_, negedge _0194_)
    if (!_0194_) _3704_ <= 6'h0c;
    else _3704_ <= { _2121_[31:29], _0356_, _0134_, _0573_ };
  assign { _1977_[25:24], _1243_, _1384_, _1669_, _0256_ } = _3704_;
  reg [64:0] _3705_;
  always_ff @(negedge _1268_, posedge _0112_)
    if (_0112_) _3705_ <= 65'h00000000000000000;
    else _3705_ <= { _0919_, _1891_[12:5], _2144_[55], _1250_, _2072_[44], _1973_[25:24], _0504_, _1597_, _0684_, _1973_[20:19], _1970_[51:20], _1253_, _1970_[18:16], _1210_, _1682_, _1970_[13:11], _2144_[4:0] };
  assign { _2280_[64:59], _1482_, _2280_[57:31], _0903_, _2280_[29:0] } = _3705_;
  reg [82:0] _3706_;
  always_ff @(negedge _1464_, negedge _0811_)
    if (!_0811_) _3706_ <= 83'h000000000000000000000;
    else _3706_ <= { _2183_[86:50], _1349_, _2183_[48:29], _2079_[21:5], _0247_, _1381_, _0241_, _1810_, _0123_, _1932_[6], _0595_, _0565_ };
  assign { _2281_[82:65], _1280_, _2281_[63:56], _1583_, _2281_[54:51], _2163_[42:25], _2281_[32:0] } = _3706_;
  reg [13:0] _3707_;
  always_ff @(posedge _0149_, posedge _0490_)
    if (_0490_) _3707_ <= 14'h22a5;
    else _3707_ <= { _2014_[12:10], _1988_[54:51], _0291_, _1988_[49], _1383_, _1988_[47:46], _1697_, _1988_[44] };
  assign { _1964_[67], _0364_, _1888_[13], _0036_, _0706_, _1888_[10:5], _0673_, _1964_[55], _1679_ } = _3707_;
  reg [25:0] _3708_;
  always_ff @(negedge _0343_, negedge _0183_)
    if (!_0183_) _3708_ <= 26'h1c1fb99;
    else _3708_ <= _1968_[44:19];
  assign { _2094_[28:26], _1779_, _2094_[24], _0691_, _1416_, _1781_, _2094_[20:19], _0545_, _2094_[17:14], _0346_, _2094_[12:6], _1767_, _2094_[4:3] } = _3708_;
  reg [7:0] _3709_;
  always_ff @(negedge _0194_, negedge _0270_)
    if (!_0270_) _3709_ <= 8'h69;
    else _3709_ <= { _0909_, _0519_, _0164_, _0635_, _0251_, _0149_, _0158_, _0207_ };
  assign _1946_[8:1] = _3709_;
  reg [11:0] _3710_;
  always_ff @(posedge _0265_, posedge _2266_[0])
    if (_2266_[0]) _3710_ <= 12'ha6a;
    else _3710_ <= { _2054_[13:9], _2254_[18], _1717_, _2254_[16:14], _1404_, _2254_[12] };
  assign { _1952_[15:12], _1385_, _1952_[10:7], _1118_, _1952_[5:4] } = _3710_;
  reg [119:0] _3711_;
  always_ff @(negedge _2021_[1], posedge _0191_)
    if (_0191_) _3711_ <= 120'h000000000000000000000000000000;
    else _3711_ <= { _2026_[11], _1097_, _2026_[9:8], _1836_, _2229_[25], _0287_, _0057_, _0665_, _2033_[23:22], _1783_, _2033_[20:6], _1407_, _2033_[4:0], _0102_, _1211_, _2281_[82:65], _1280_, _2281_[63:56], _1583_, _2281_[54:51], _2163_[42:25], _2281_[32:0], _0046_, _1235_ };
  assign { _2282_[119:102], _0938_, _2282_[100:99], _2160_[50:24], _2282_[71:60], _2149_[60:20], _2282_[18:11], _1444_, _2282_[9:0] } = _3711_;
  reg [102:0] _3712_;
  always_ff @(negedge _0217_, negedge _0379_)
    if (!_0379_) _3712_ <= 103'h00000000000000000000000000;
    else _3712_ <= { _1901_[72:70], _1978_[13:7], _0277_, _0096_, _0184_, _2019_[58:57], _1636_, _2019_[55:37], _0070_, _1920_[31:22], _0056_, _1920_[20:19], _1816_, _1920_[17:16], _1168_, _1920_[14:2], _2019_[5], _1942_[86:58], _1006_, _1077_, _0248_, _1684_, _2028_[3], _1326_, _2028_[1] };
  assign { _2102_[115:53], _0399_, _2102_[51:34], _1662_, _2102_[32:13] } = _3712_;
  reg [20:0] _3713_;
  always_ff @(posedge _0607_, posedge _0113_)
    if (_0113_) _3713_ <= 21'h08f66f;
    else _3713_ <= { _2102_[86:70], _0306_, _0620_, _0686_, _0151_ };
  assign { _2221_[76:75], _0536_, _2221_[73:71], _1688_, _1815_, _1432_, _2221_[67:59], _1543_, _2221_[57:56] } = _3713_;
  reg [21:0] _3714_;
  always_ff @(posedge _1017_, negedge _1888_[9])
    if (!_1888_[9]) _3714_ <= 22'h1f63ae;
    else _3714_ <= { _2101_[34], _0005_, _1205_, _0116_, _0386_, _0192_, _0157_, _0196_, _2003_[10:9], _1126_, _1631_, _2003_[6:3], _1372_, _1217_, _2003_[0], _0286_, _0640_, _0672_ };
  assign { _2151_[25], _2146_[23:21], _1763_, _2146_[19:4], _2151_[4] } = _3714_;
  reg [14:0] _3715_;
  always_ff @(posedge _0102_, negedge _0084_)
    if (!_0084_) _3715_ <= 15'h6c0c;
    else _3715_ <= { _2054_[33:31], _1683_, _2054_[29], _0561_, _1530_, _0588_, _1890_[11], _0350_, _0716_, _1890_[8:6], _0294_ };
  assign { _1601_, _2107_[14:13], _2092_[14:7], _1548_, _2092_[5], _2107_[2:1] } = _3715_;
  always_ff @(negedge _0317_, posedge _1464_)
    if (_1464_) _1470_ <= 1'h1;
    else _1470_ <= _1550_;
  reg [120:0] _3717_;
  always_ff @(posedge _1634_, posedge _0159_)
    if (_0159_) _3717_ <= 121'h0000000000000000000000000000000;
    else _3717_ <= { _0133_, _0283_, _0566_, _1994_[9:6], _0840_, _1994_[4:3], _0597_, _2048_[51:50], _1423_, _2048_[48:47], _2005_[10:8], _1327_, _2005_[6:4], _2048_[39:38], _1150_, _2048_[36], _1010_, _2048_[34:17], _1368_, _1627_, _0919_, _0811_, _0193_, _1470_, _0730_, _0669_, _0211_, _1518_, _0436_, _0241_, _0283_, _2065_[57:40], _1400_, _2065_[38:27], _1430_, _2065_[25:0], _0039_, _0238_, _0269_, _0076_ };
  assign { _2283_[120:86], _1240_, _2283_[84:70], _2129_, _2283_[52:18], _0365_, _2283_[16:0] } = _3717_;
  reg [12:0] _3718_;
  always_ff @(negedge _0656_, posedge out_data[1344])
    if (out_data[1344]) _3718_ <= 13'h0bc0;
    else _3718_ <= { _2033_[11:8], _0675_, _0152_, _1956_[18:15], _0506_, _1956_[13:12] };
  assign { _1901_[15:14], _0760_, _1901_[12:10], _0879_, _1901_[8:5], _1078_, _1901_[3] } = _3718_;
  reg [40:0] _3719_;
  always_ff @(negedge _2112_[90], posedge _0069_)
    if (_0069_) _3719_ <= 41'h000750b17a3;
    else _3719_ <= { _1981_[11:9], _0299_, _0223_, _1981_[6:4], _1589_, _1096_, _0247_, _1980_[23:6], _1367_, _1980_[4], _1681_, _1980_[2:0], _1003_, _0207_, _0164_, _0317_, _0219_, _1174_ };
  assign { _2284_[40], _1477_, _2284_[38:32], _1143_, _2284_[30:7], _1437_, _2284_[5:0] } = _3719_;
  reg [81:0] _3720_;
  always_ff @(posedge _1970_[50], negedge _1575_)
    if (!_1575_) _3720_ <= 82'h000000000000000000000;
    else _3720_ <= { _2094_[130:103], _1291_, _2094_[101:94], _1263_, _2094_[92:69], _0361_, _1130_, _0038_, _0033_, _2275_, _0185_, _1551_ };
  assign { _2285_[81:76], _1398_, _2285_[74:71], _1611_, _2285_[69:55], _2248_[35:7], _2285_[25:0] } = _3720_;
  reg [6:0] _3721_;
  always_ff @(posedge _0907_, posedge _1900_[82])
    if (_1900_[82]) _3721_ <= 7'h7d;
    else _3721_ <= { _1888_[10:6], _1013_, _0873_ };
  assign { _2145_[7], _1062_, _2145_[5], _1635_, _2145_[3:1] } = _3721_;
  reg [14:0] _3722_;
  always_ff @(negedge _0082_, posedge _1561_)
    if (_1561_) _3722_ <= 15'h5f8a;
    else _3722_ <= { _0219_, _0685_, _0289_, _2061_[10:4], _1554_, _2061_[2:0], _0351_ };
  assign { _2286_[14:9], _0966_, _2286_[7:6], _1146_, _2286_[4:0] } = _3722_;
  reg [99:0] _3723_;
  always_ff @(negedge _0228_, posedge _0733_)
    if (_0733_) _3723_ <= 100'h0000000000000000000000000;
    else _3723_ <= { _2112_[89:81], _2095_[130:127], _2007_[8:1], _1441_, _2095_[117:116], _1046_, _0025_, _0189_, _0316_, _0043_, _0226_, _0096_, _0022_, _0237_, _0125_, _0125_, _0356_, _0152_, _0200_, _0227_, _0068_, _0152_, _0043_, _0103_, _0043_, _0043_, _0265_, _0134_, _0189_, _0103_, _0316_, _0463_, _0125_, _0134_, _0490_, _0033_, _0918_, _0463_, _0106_, _0265_, _1964_[67], _0364_, _1888_[13], _0036_, _0706_, _1888_[10:5], _0673_, _1964_[55], _1679_, _0226_, _0200_, _0926_, _0674_, _0610_, _2067_[2:1], _0775_, _0316_, _0287_, _0043_, _0191_, _0103_, _0132_, _0068_, _0128_, _0128_, _0356_, _0733_, _0277_, _0356_, _0134_, _0189_, _0096_, _0221_, _0316_, _1283_ };
  assign { _2216_[100:99], _1511_, _2216_[97:86], _0734_, _2216_[84:80], _1278_, _2216_[78:62], _1952_[215:214], _1083_, _1952_[212:206], _1246_, _1952_[204:184], _1389_, _1952_[182:177], _0344_, _1952_[175:165], _1194_, _1952_[163:157], _2216_[2:1] } = _3723_;
  reg [29:0] _3724_;
  always_ff @(posedge _0450_, posedge _2146_[19])
    if (_2146_[19]) _3724_ <= 30'h00b9853a;
    else _3724_ <= { _2216_[83:80], _1278_, _2216_[78:62], _1952_[215:214], _1083_, _1952_[212:209], _0178_ };
  assign { _2287_[29:26], _0500_, _2287_[24:23], _0720_, _2287_[21:16], _2180_, _2287_[8:0] } = _3724_;
  reg [1:0] _3725_;
  always_ff @(posedge _0151_, negedge _0206_)
    if (!_0206_) _3725_ <= 2'h1;
    else _3725_ <= { _0113_, _0025_ };
  assign _2126_[44:43] = _3725_;
  reg [5:0] _3726_;
  always_ff @(negedge _1347_, negedge _0152_)
    if (!_0152_) _3726_ <= 6'h35;
    else _3726_ <= { _1812_, _1675_, _0287_, _0586_, _0634_, _0103_ };
  assign { _1951_[123], _1122_, _1951_[121:119], _1609_ } = _3726_;
  reg [21:0] _3727_;
  always_ff @(posedge _0946_, posedge _2030_[13])
    if (_2030_[13]) _3727_ <= 22'h26df18;
    else _3727_ <= { _2032_[18:13], _0606_, _2032_[11:10], _0420_, _0649_, _0651_, _0692_, _0317_, _1009_, _0587_, _0489_, _1046_, _0102_, _0211_, _1283_, _0678_ };
  assign { _1943_[81:75], _1082_, _1943_[73:68], _1504_, _1943_[66:64], _1724_, _1943_[62:60] } = _3727_;
  reg [4:0] _3728_;
  always_ff @(negedge _0997_, posedge _0988_)
    if (_0988_) _3728_ <= 5'h0c;
    else _3728_ <= { _0652_, _0873_, _1114_, _0999_, _0808_ };
  assign { _2288_[4], _0491_, _2288_[2], _1622_, _2288_[0] } = _3728_;
  reg [14:0] _3729_;
  always_ff @(negedge _1047_, negedge _0220_)
    if (!_0220_) _3729_ <= 15'h6e17;
    else _3729_ <= { _2121_[25:22], _2031_[66], _0328_, _2031_[64], _0007_, _1699_, _2031_[61:58], _0096_, _0038_ };
  assign _1964_[21:7] = _3729_;
  reg [16:0] _3730_;
  always_ff @(negedge _1311_, posedge _1064_)
    if (_1064_) _3730_ <= 17'h0d2e4;
    else _3730_ <= { in_data[96:81], _0194_ };
  assign { _2120_[32:30], _1762_, _2120_[28:16] } = _3730_;
  reg [121:0] _3731_;
  always_ff @(negedge _1345_, negedge _1047_)
    if (!_1047_) _3731_ <= 122'h0000000000000000000000000000000;
    else _3731_ <= { _1980_[9:6], _1367_, _1645_, _0165_, _0099_, _0096_, _0489_, _1374_, _0993_, _0403_, _2017_[65:61], _1364_, _2017_[59:37], _1410_, _2017_[35:33], _0414_, _2017_[31:14], _1442_, _2017_[12:0], _0841_, _0222_, _0448_, _1205_, _2139_[49], _1748_, _2139_[47:45], _1837_, _2139_[43], _1256_, _2139_[41:40], _2046_[6], _1756_, _2046_[4], _1094_, _2046_[2:0], _0946_, _0186_, _1909_[12], _1908_[39:38], _1885_, _1908_[36], _1270_, _1908_[34], _1048_, _1909_[4:2], _1167_, _0550_, _0709_, _0918_, _0175_, _0218_, _1561_, _0816_, _0220_ };
  assign { _2289_[121], _2143_[84:77], _1759_, _2143_[75:3], _2150_[26:0], _2289_[11:0] } = _3731_;
  reg [8:0] _3732_;
  always_ff @(posedge _0132_, negedge _0232_)
    if (!_0232_) _3732_ <= 9'h043;
    else _3732_ <= { _2170_[82:80], _1977_[25:24], _1243_, _1384_, _1669_, _0256_ };
  assign { _1530_, _0588_, _1890_[11], _0350_, _0716_, _1890_[8:6], _0294_ } = _3732_;
  reg [10:0] _3733_;
  always_ff @(negedge _0343_, negedge _0182_)
    if (!_0182_) _3733_ <= 11'h768;
    else _3733_ <= { _1955_[24:21], _0325_, _0053_, _0161_, _0385_, _0919_, _1518_, _0348_ };
  assign { _2094_[55:47], _1732_, _2094_[45] } = _3733_;
  reg [60:0] _3734_;
  always_ff @(negedge _0625_, negedge _1175_)
    if (!_1175_) _3734_ <= 61'h1ffffffffc6e35e9;
    else _3734_ <= { _2064_[19:14], _1004_, _0746_, _0132_, _0132_, _0187_, _1322_, _1247_, _0082_, _1951_[123], _1122_, _1951_[121:119], _1609_, _0048_, _0611_, _0481_, _2288_[4], _0491_, _2288_[2], _1622_, _2288_[0], _0438_, _1527_, _0270_, _2088_[22:20], _0577_, _2088_[18:0], _1956_[18:15], _0506_, _1956_[13:12] };
  assign { _2095_[86:40], _1516_, _2095_[38:26] } = _3734_;
  reg [14:0] _3735_;
  always_ff @(negedge _0656_, negedge _0695_)
    if (!_0695_) _3735_ <= 15'h4274;
    else _3735_ <= { _1323_, _2001_[109], _1309_, _1081_, _2001_[106:103], _1351_, _2001_[101:99], _0134_, _1405_, _0024_ };
  assign { _2236_[39:32], _1700_, _2236_[30:25] } = _3735_;
  reg [17:0] _3736_;
  always_ff @(posedge _0266_, negedge _1247_)
    if (!_1247_) _3736_ <= 18'h19ad1;
    else _3736_ <= { _1911_[14:8], _1284_, _0908_, _2063_[28], _2081_[21], _1269_, _2081_[19], _0905_, _0632_, _1266_, _0887_, _0991_ };
  assign { _2108_[32:31], _1414_, _2108_[29:15] } = _3736_;
  reg [52:0] _3737_;
  always_ff @(negedge _0661_, posedge _0611_)
    if (_0611_) _3737_ <= 53'h1fffffb22c59d1;
    else _3737_ <= { _1979_[40:22], _0790_, _0146_, _0730_, _0134_, _0105_, _1964_[52], _1795_, _1964_[50:48], _1016_, _1964_[46:45], _0492_, _1964_[43], _1706_, _0306_, _1114_, _1066_, _0915_, _0613_, _1808_, _0099_, _0198_, _1936_[47:44], _1612_, _1936_[42], _0418_, _1936_[40], _0268_, _0781_ };
  assign { _2290_[52:46], _2097_[39:5], _2290_[10:0] } = _3737_;
  reg [23:0] _3738_;
  always_ff @(posedge _0176_, negedge _1951_[168])
    if (!_1951_[168]) _3738_ <= 24'h6cab26;
    else _3738_ <= { _1975_[54], _1790_, _1339_, _1836_, _2229_[25], _0704_, _1402_, _0216_, _0694_, _0209_, _0518_, _1750_, _2003_[10:9], _1126_, _1631_, _2003_[6:3], _1372_, _1217_, _2003_[0], _0540_ };
  assign { _2291_[23:11], _1628_, _2291_[9:0] } = _3738_;
  reg [1:0] _3739_;
  always_ff @(negedge _0149_, negedge _2269_[12])
    if (!_2269_[12]) _3739_ <= 2'h0;
    else _3739_ <= { _0724_, _0140_ };
  assign { _1709_, _2292_[0] } = _3739_;
  reg [38:0] _3740_;
  always_ff @(negedge _0715_, negedge _1390_)
    if (!_1390_) _3740_ <= 39'h7f9fb93cbc;
    else _3740_ <= { _1994_[3], _0597_, _2048_[51:50], _1423_, _2048_[48:47], _2005_[10:8], _1327_, _2005_[6:4], _2048_[39:38], _1150_, _2048_[36], _1010_, _2048_[34:18], _0801_, _0214_, _0134_ };
  assign { _2101_[93:90], _0910_, _2101_[88], _1895_[35:26], _1111_, _1895_[24:20], _1757_, _1895_[18:3] } = _3740_;
  reg [14:0] _3741_;
  always_ff @(negedge _0648_, posedge _1322_)
    if (_1322_) _3741_ <= 15'h1111;
    else _3741_ <= { _2261_[89:78], _1396_, _1131_, _0251_ };
  assign { _2293_[14:13], _2166_[46], _1100_, _2166_[44:36], _2293_[1:0] } = _3741_;
  reg [1:0] _3742_;
  always_ff @(posedge _0019_, posedge _0401_)
    if (_0401_) _3742_ <= 2'h3;
    else _3742_ <= { _0672_, _0799_ };
  assign { _0844_, _1713_ } = _3742_;
  reg [13:0] _3743_;
  always_ff @(posedge _2015_[17], negedge _1561_)
    if (!_1561_) _3743_ <= 14'h152b;
    else _3743_ <= { _0335_, _0510_, _0692_, _0272_, _0613_, _0189_, _0298_, _0941_, _1716_, _1996_[4], _1365_, _0104_, _1476_, _1467_ };
  assign { _2294_[13:6], _0520_, _2294_[4], _1140_, _2294_[2:0] } = _3743_;
  reg [31:0] _3744_;
  always_ff @(posedge _0891_, negedge _1345_)
    if (!_1345_) _3744_ <= 32'd787237412;
    else _3744_ <= { _2134_[4:3], _2194_[4], _1091_, _2205_[9:3], _0718_, _1343_, _0919_, _2108_[32:31], _1414_, _2108_[29:15] };
  assign { _2237_[31:29], _1219_, _2237_[27:0] } = _3744_;
  reg [31:0] _3745_;
  always_ff @(posedge _1247_, negedge _1976_[2])
    if (!_1976_[2]) _3745_ <= 32'd923118282;
    else _3745_ <= { _2080_[30:23], _0008_, _2080_[21:12], _0325_, _0214_, _0726_, _0138_, _0988_, _1061_, out_data[896], _1390_, _0328_, _0289_, _0666_, _1470_, _0080_ };
  assign { _2295_[31:28], _0002_, _2295_[26:12], _0750_, _2295_[10:0] } = _3745_;
  reg [8:0] _3746_;
  always_ff @(negedge _1991_[53], posedge _1972_[20])
    if (_1972_[20]) _3746_ <= 9'h1bd;
    else _3746_ <= { _1053_, _0032_, _1055_, _0625_, _0386_, _1283_, _0419_, _0801_, _0270_ };
  assign { _2117_[8:6], _0432_, _2117_[4:1], _2213_[3] } = _3746_;
  reg [43:0] _3747_;
  always_ff @(negedge _0101_, negedge _0241_)
    if (!_0241_) _3747_ <= 44'h0001ac52f25;
    else _3747_ <= { in_data[1102:1072], _0025_, _0189_, _0101_, _0189_, _0025_, _1716_, _1996_[4], _1365_, _0104_, _1476_, _1467_, _0200_, _0101_ };
  assign { _2121_[43:39], _0864_, _1346_, _2121_[36:35], _1600_, _2121_[33:28], _0653_, _2121_[26:22], _2031_[66], _0328_, _2031_[64], _0007_, _1699_, _2031_[61:55], _1806_, _2031_[53], _0206_, _2031_[51], _1800_, _2031_[49:47], _2121_[1:0] } = _3747_;
  reg [31:0] _3748_;
  always_ff @(negedge _0287_, negedge _1000_)
    if (!_1000_) _3748_ <= 32'd3481360913;
    else _3748_ <= { _0237_, _0227_, _0127_, _0304_, _0320_, _0097_, _0573_, _0317_, _0197_, _1716_, _1996_[4], _1365_, _0104_, _1476_, _1467_, _0690_, _0237_, _0189_, _0194_, _0106_, _0287_, _1254_, _0468_, _2006_[6], _0404_, _2006_[4:3], _1931_[3], _1308_, _0513_, _0082_, _0306_ };
  assign { _2063_[43], _1615_, _0147_, _2063_[40:38], _1911_[14:8], _1284_, _0908_, _2063_[28], _2081_[21], _1269_, _2081_[19], _1376_, _2081_[17:16], _0642_, _2240_[9:1] } = _3748_;
  reg [4:0] _3749_;
  always_ff @(negedge _2006_[6], posedge _0661_)
    if (_0661_) _3749_ <= 5'h0e;
    else _3749_ <= { _1441_, _2095_[117:114] };
  assign { _1786_, _0402_, _1397_, _1569_, _1970_[5] } = _3749_;
  reg [7:0] _3750_;
  always_ff @(posedge _0116_, posedge _1901_[8])
    if (_1901_[8]) _3750_ <= 8'hcc;
    else _3750_ <= { _2048_[50], _0537_, _0228_, _0642_, _0605_, _0312_, _1609_, _0212_ };
  assign { _2149_[13:8], _1152_, _2149_[6] } = _3750_;
  reg [19:0] _3751_;
  always_ff @(negedge _0191_, negedge _0690_)
    if (!_0690_) _3751_ <= 20'hdd489;
    else _3751_ <= { _2001_[111], _1323_, _2001_[109], _1309_, _1081_, _2001_[106:103], _1351_, _2001_[101:99], _1353_, _2001_[97], _1359_, _0277_, _0134_, _0043_, _0150_ };
  assign { _2205_[19:18], _0726_, _2194_[9], _2134_[6], _0003_, _2134_[4:3], _2194_[4], _1091_, _2205_[9:3], _1693_, _2205_[1:0] } = _3751_;
  reg [10:0] _3752_;
  always_ff @(posedge _1130_, negedge _2094_[111])
    if (!_2094_[111]) _3752_ <= 11'h6d7;
    else _3752_ <= { _1153_, _1893_[10:7], _1034_, _1893_[5:4], _1374_, _1787_, _0126_ };
  assign { _2296_[10:7], _1581_, _2296_[5:4], _0388_, _2296_[2:0] } = _3752_;
  reg [1:0] _3753_;
  always_ff @(posedge _0469_, posedge _1025_)
    if (_1025_) _3753_ <= 2'h2;
    else _3753_ <= _1951_[129:128];
  assign { _2165_[11], _1187_ } = _3753_;
  reg [14:0] _3754_;
  always_ff @(posedge _0525_, posedge _0296_)
    if (_0296_) _3754_ <= 15'h0f04;
    else _3754_ <= { _0311_, _0986_, _1908_[14:13], _1564_, _1908_[11:10], _0535_, _1908_[8:7], _1818_, _0727_, _1231_, _0071_, _0116_ };
  assign { _1927_[19], _1565_, _1927_[17:6], _0853_ } = _3754_;
  reg [24:0] _3755_;
  always_ff @(negedge _0325_, posedge _1464_)
    if (_1464_) _3755_ <= 25'h06d4425;
    else _3755_ <= { _1959_[7], _1202_, _0899_, _0793_, _2221_[76:75], _0536_, _2221_[73:71], _1688_, _1815_, _1432_, _2221_[67:59], _1543_, _2221_[57:56] };
  assign { _2297_[24:3], _1735_, _2297_[1:0] } = _3755_;
  reg [29:0] _3756_;
  always_ff @(posedge _1913_[11], posedge _0295_)
    if (_0295_) _3756_ <= 30'h211b3de4;
    else _3756_ <= { _2021_[16:13], _1189_, _2021_[11:6], _1405_, _0166_, _2286_[14:9], _0966_, _2286_[7:6], _1146_, _2286_[4:0], _0096_, _1585_ };
  assign { _1954_[28:12], _1872_, _1954_[10:9], out_data[1952], _1954_[7:0], _2298_[0] } = _3756_;
  reg [26:0] _3757_;
  always_ff @(posedge _0026_, negedge _1345_)
    if (!_1345_) _3757_ <= 27'h24c52b5;
    else _3757_ <= { _2058_[79:60], _1427_, _2058_[58:54], _0353_ };
  assign { _2299_[26:9], _1271_, _2299_[7:0] } = _3757_;
  reg [4:0] _3758_;
  always_ff @(negedge _0134_, negedge _0067_)
    if (!_0067_) _3758_ <= 5'h0d;
    else _3758_ <= { _0119_, _1038_, _0182_, _0108_, _0999_ };
  assign _1915_[10:6] = _3758_;
  reg [25:0] _3759_;
  always_ff @(negedge _0103_, negedge _0025_)
    if (!_0025_) _3759_ <= 26'h285ee6c;
    else _3759_ <= { _2287_[29:26], _0500_, _2287_[24:23], _0720_, _2287_[21:16], _2180_, _2287_[8:5], _1310_ };
  assign _2139_[26:1] = _3759_;
  reg [21:0] _3760_;
  always_ff @(posedge _0202_, negedge _2001_[126])
    if (!_2001_[126]) _3760_ <= 22'h12b37e;
    else _3760_ <= { _2121_[22], _2031_[66], _0328_, _2031_[64], _0007_, _1699_, _2031_[61:55], _1806_, _2031_[53], _0206_, _2031_[51], _1800_, _2031_[49:47], _2121_[1] };
  assign { _2227_[22:12], _2211_[13:7], _1541_, _2211_[5:3] } = _3760_;
  reg [24:0] _3761_;
  always_ff @(negedge _0345_, posedge _1980_[17])
    if (_1980_[17]) _3761_ <= 25'h17850a0;
    else _3761_ <= { _2138_[62:39], _0773_ };
  assign { _2300_[24:15], _1730_, _2300_[13:0] } = _3761_;
  reg [9:0] _3762_;
  always_ff @(negedge _1377_, negedge _1056_)
    if (!_1056_) _3762_ <= 10'h1e7;
    else _3762_ <= { _2149_[57:50], _0766_, _0631_ };
  assign { _2197_[91:90], _0877_, _2197_[88:82] } = _3762_;
  reg [24:0] _3763_;
  always_ff @(posedge _0873_, negedge _0678_)
    if (!_0678_) _3763_ <= 25'h15b1e77;
    else _3763_ <= { _2132_[1], _0791_, _2258_[14:0], _0967_, _0354_, _2126_[44:43], _0578_, _1067_, _0993_, _0403_ };
  assign { _2301_[24:23], _2173_[23:21], _1460_, _2173_[19:3], _2301_[1:0] } = _3763_;
  reg [55:0] _3764_;
  always_ff @(posedge _0455_, posedge _0152_)
    if (_0152_) _3764_ <= 56'h00000012058fce;
    else _3764_ <= { _0038_, _2139_[35:32], _1354_, _1054_, _2139_[29:27], _2103_, _1651_, _0292_, _1043_, _0598_, _0185_, _1130_, _1084_, _1422_, _0675_, _0215_, _0164_, _1799_, _0277_, _0531_, _1000_, _0531_, _1076_, _1639_, _1900_[46:37], _0767_, _1900_[35:29], _0230_, _1833_, _1900_[26] };
  assign { _2302_[55:53], _2159_[50:48], _1907_[55:25], _1535_, _1907_[23:16], _2159_[7:2], _1842_, _2159_[0], _2302_[1:0] } = _3764_;
  reg [15:0] _3765_;
  always_ff @(negedge _0018_, negedge _0993_)
    if (!_0993_) _3765_ <= 16'had65;
    else _3765_ <= { _1987_[32:31], _0693_, _1987_[29:23], _0798_, _1987_[21:19], _1835_, _0113_ };
  assign { _1898_[15:10], _0765_, _1898_[8:0] } = _3765_;
  reg [5:0] _3766_;
  always_ff @(posedge _0599_, posedge _0749_)
    if (_0749_) _3766_ <= 6'h06;
    else _3766_ <= { _0635_, _1027_, _0065_, _0987_, _0656_, _0132_ };
  assign { _0063_, _2232_[6:5], _0375_, _2232_[3], _1544_ } = _3766_;
  reg [11:0] _3767_;
  always_ff @(negedge _0671_, posedge _1561_)
    if (_1561_) _3767_ <= 12'h6a1;
    else _3767_ <= { _2291_[20:11], _1628_, _2291_[9] };
  assign { _1887_[11:10], _1850_, _1887_[8], _1537_, _1887_[6:0] } = _3767_;
  reg [60:0] _3768_;
  always_ff @(posedge _0028_, posedge _0408_)
    if (_0408_) _3768_ <= 61'h1ffffffffccb8119;
    else _3768_ <= { _2165_[11], _0816_, _0157_, _1831_, _0166_, _1424_, _1399_, _2262_[56:54], _1690_, _2262_[52], _2025_[43:40], _1785_, _2025_[38:34], _1510_, _2025_[32:27], _0896_, _2025_[25], _1556_, _0114_, _0319_, _2041_[32:31], _1755_, _2041_[29:24], _0233_, _0499_, _2114_[25:23], _0633_, _0162_, _1959_[7], _1202_, _0918_, _0229_, _1935_[18:17], _0558_, _1935_[15], out_data[1344], _0321_, _0175_ };
  assign { _2303_[60:7], _1859_, _2303_[5:0] } = _3768_;
  reg [33:0] _3769_;
  always_ff @(posedge _1211_, posedge _0177_)
    if (_0177_) _3769_ <= 34'h05bda4628;
    else _3769_ <= { _1309_, _1081_, _2001_[106:103], _1351_, _0194_, _0121_, _0096_, _0228_, _0227_, _2000_[20:19], _0564_, _2000_[17:14], _0925_, _1939_[12:8], _0501_, _1939_[6], _1306_, _2000_[4:3], _1632_, _1373_, _2000_[0], _0311_ };
  assign { _2000_[59:50], _1570_, _2000_[48:46], _1314_, _1419_, _0391_, _2000_[42:35], _1747_, _2000_[33:31], _1307_, _2000_[29:27], _1318_ } = _3769_;
  reg [24:0] _3770_;
  always_ff @(posedge _0659_, posedge _0670_)
    if (_0670_) _3770_ <= 25'h1a35f5f;
    else _3770_ <= { _2053_[31:28], _1667_, _0297_, _0784_, _1015_, _1144_, _1084_, _1179_, _1051_, _0238_, _1044_, _0276_, _0561_, _0150_, _0636_, _0709_, out_data[1184], _0186_, _1409_, _0012_, _0337_, _0027_ };
  assign { _1942_[47:45], _1285_, _1942_[43:39], _1547_, _1942_[37:23] } = _3770_;
  always_ff @(posedge _0871_, posedge _0565_)
    if (_0565_) _2304_ <= 3'h1;
    else _2304_ <= { _0134_, _0095_, _0637_ };
  reg [26:0] _3772_;
  always_ff @(posedge _1746_, posedge _0475_)
    if (_0475_) _3772_ <= 27'h39845da;
    else _3772_ <= { _2064_[35:34], _2024_[13:12], _1825_, _2024_[10:2], _2064_[21:14], _1676_, _2064_[12], _1951_[130:128] };
  assign { _2251_[16:15], _1490_, _2214_[22], _2251_[12:1], _2305_[10:0] } = _3772_;
  reg [43:0] _3773_;
  always_ff @(posedge _0091_, posedge _0898_)
    if (_0898_) _3773_ <= 44'h0005d73a399;
    else _3773_ <= { _0726_, _2108_[32:31], _1414_, _2108_[29:15], _0318_, _1422_, _1549_, _2117_[8:6], _0432_, _2117_[4:1], _2213_[3], _0269_, _0425_, _1722_, _0018_, _0180_, _0646_, _1077_, _0248_, _1684_, _2028_[3], _1326_, _2028_[1], _1551_ };
  assign { _2306_[43:26], _1854_, _2306_[24:0] } = _3773_;
  reg [29:0] _3774_;
  always_ff @(negedge _0094_, negedge _0489_)
    if (!_0489_) _3774_ <= 30'h1b0f447b;
    else _3774_ <= { _2080_[23], _0008_, _2080_[21:15], _0745_, _2022_[8:6], _1160_, _2022_[4:3], _1069_, _2022_[1:0], _1046_, _1245_, _0044_, _0152_, _0351_, _0134_, _0220_, _0228_, _0022_, _1362_, _0115_ };
  assign { _2307_[29:24], _1576_, _2307_[22], _0428_, _2307_[20:10], _1856_, _2307_[8:0] } = _3774_;
  reg [10:0] _3775_;
  always_ff @(posedge _0134_, posedge _1922_[1])
    if (_1922_[1]) _3775_ <= 11'h792;
    else _3775_ <= { _1600_, _2121_[33:28], _0653_, _2121_[26], _1046_, _0227_ };
  assign { _1981_[11:9], _0299_, _0223_, _1981_[6:2], _1794_ } = _3775_;
  reg [11:0] _3776_;
  always_ff @(negedge _1465_, posedge _1663_)
    if (_1663_) _3776_ <= 12'h70c;
    else _3776_ <= { _1907_[28:25], _1535_, _1907_[23:17] };
  assign _2161_[11:0] = _3776_;
  reg [17:0] _3777_;
  always_ff @(negedge _1942_[8], posedge _0919_)
    if (_0919_) _3777_ <= 18'h1e1a8;
    else _3777_ <= { _2294_[13:6], _0520_, _2294_[4], _1140_, _1552_, _0475_, _0324_, _0228_, _1484_, _1770_, _1935_[47] };
  assign { _2177_[17:15], _1495_, _2177_[13:5], _1191_, _2177_[3:0] } = _3777_;
  reg [9:0] _3778_;
  always_ff @(negedge _0242_, posedge _1136_)
    if (_1136_) _3778_ <= 10'h0b5;
    else _3778_ <= { _1889_[2:1], _1363_, _0000_, _1134_, _0481_, _0905_, _0411_, _0221_, _0936_ };
  assign { _2183_[12:9], _0906_, _2183_[7:3] } = _3778_;
  reg [1:0] _3779_;
  always_ff @(posedge _0717_, negedge _1956_[15])
    if (!_1956_[15]) _3779_ <= 2'h2;
    else _3779_ <= { _1891_[7], _0032_ };
  assign { _1916_[6], _1656_ } = _3779_;
  reg [23:0] _3780_;
  always_ff @(posedge _0578_, posedge _0713_)
    if (_0713_) _3780_ <= 24'hd2a69e;
    else _3780_ <= { _1984_[36], _0251_, _1984_[34:31], _0591_, _0772_, _0438_, _0176_, _1112_, out_data[896], _0318_, _1102_, _1377_, _0315_, _1108_, _2089_[5:4], _1769_, _2089_[2], _1526_, _0011_, _0306_ };
  assign { _2178_[42:26], _0396_, _2178_[24:19] } = _3780_;
  reg [49:0] _3781_;
  always_ff @(negedge _0984_, posedge _0232_)
    if (_0232_) _3781_ <= 50'h00000612e3754;
    else _3781_ <= { _2281_[73:65], _1280_, _2281_[63:56], _1583_, _2281_[54:51], _2163_[42:25], _2281_[32], _0116_, _0071_, _1424_, _1096_, _1549_, _0193_, _1655_, _0799_ };
  assign { _2231_[94:81], _2200_[47:42], _1855_, _0923_, _2200_[39:20], _2231_[52:45] } = _3781_;
  reg [51:0] _3782_;
  always_ff @(negedge _1472_, negedge _0018_)
    if (!_0018_) _3782_ <= 52'h0000045e80581;
    else _3782_ <= { _2271_[11:6], _0374_, _1671_, _2203_[16:10], _1571_, _2203_[8], _1938_[8:5], _0131_, _2203_[2:0], _0866_, _1841_, _0652_, _0751_, _1435_, _0203_, _0416_, _0792_, _0306_, _0067_, _0746_, _0195_, _0272_, _1598_, _0058_, _2304_, _0342_, _0458_, _0338_, _0561_, _0689_, _0208_, _0216_, _0994_, _0756_ };
  assign _2197_[77:26] = _3782_;
  reg [104:0] _3783_;
  always_ff @(negedge _1063_, negedge _1708_)
    if (!_1708_) _3783_ <= 105'h000000000000000000000000000;
    else _3783_ <= { _2270_[69:67], _0667_, _2094_[130:103], _1291_, _2094_[101:94], _1263_, _2094_[92:73], _1675_, _1429_, _0112_, _0022_, _0490_, _0152_, _0043_, _0032_, _1451_, _1065_, _0250_, _2299_[26:9], _1271_, _2299_[7:0], _1298_, _0714_, _0663_, _0662_, _0454_ };
  assign { _2308_[104:100], _2178_[81:79], _1903_[38:36], _1213_, _1903_[34:3], _2308_[60:0] } = _3783_;
  reg [7:0] _3784_;
  always_ff @(negedge _1081_, posedge _0153_)
    if (_0153_) _3784_ <= 8'h3d;
    else _3784_ <= { _1988_[33], _0208_, _0018_, _0057_, _1076_, _0046_, _0769_, _0566_ };
  assign { _1933_[13:9], _1244_, _1933_[7:6] } = _3784_;
  reg [12:0] _3785_;
  always_ff @(posedge _2021_[9], posedge _2146_[12])
    if (_2146_[12]) _3785_ <= 13'h1451;
    else _3785_ <= { _2139_[22:16], _0353_, _0663_, _0303_, _0537_, _0254_, _0210_ };
  assign { _2309_[12:7], _1874_, _2309_[5], _1180_, _2309_[3:0] } = _3785_;
  reg [11:0] _3786_;
  always_ff @(negedge _2156_[78], negedge _1233_)
    if (!_1233_) _3786_ <= 12'h03e;
    else _3786_ <= { _1927_[15:11], _1835_, _0052_, _1935_[18:17], _0558_, _1935_[15], _1315_ };
  assign { _0471_, _2226_[33:24], _1921_ } = _3786_;
  reg [19:0] _3787_;
  always_ff @(posedge _2075_[11], posedge _0176_)
    if (_0176_) _3787_ <= 20'hf9703;
    else _3787_ <= _2153_[22:3];
  assign { _2188_[24:19], _0459_, _2188_[17:5] } = _3787_;
  reg [61:0] _3788_;
  always_ff @(posedge _0779_, posedge _0191_)
    if (_0191_) _3788_ <= 62'h0000000072016e47;
    else _3788_ <= { _1903_[23:18], _1117_, _1021_, _0529_, _0206_, _0253_, _1086_, _1339_, _0134_, _2133_[6:1], _1727_, _1129_, _0670_, _0683_, _0944_, _2172_, _1006_, _0786_, _1120_, _2044_[8:6], _0668_, _2044_[4:1], _1461_, _0640_ };
  assign { _2310_[61:50], _2195_[10:6], _2310_[44:14], _2181_[11:2], _2310_[3:0] } = _3788_;
  reg [2:0] _3789_;
  always_ff @(posedge _0816_, posedge _2140_[11])
    if (_2140_[11]) _3789_ <= 3'h1;
    else _3789_ <= { _0716_, _1392_, _0373_ };
  assign { _2186_[3:2], _0932_ } = _3789_;
  reg [1:0] _3790_;
  always_ff @(negedge _0552_, posedge _0354_)
    if (_0354_) _3790_ <= 2'h3;
    else _3790_ <= { _0166_, _1363_ };
  assign { _1914_[10], _1529_ } = _3790_;
  reg [43:0] _3791_;
  always_ff @(posedge _0082_, negedge _0638_)
    if (!_0638_) _3791_ <= 44'h0005d3dafd0;
    else _3791_ <= { _2170_[80:70], _2070_[32:18], _1201_, _2070_[16:11], _1796_, _2070_[9:5], _0165_, _2070_[3:1], _0529_ };
  assign { _1070_, _2245_[79], _1313_, _0624_, _2141_[22:19], _2245_[72:70], _1984_[46:39], _1714_, _1984_[37:36], _0251_, _1984_[34:15], _2245_[37] } = _3791_;
  reg [55:0] _3792_;
  always_ff @(negedge _1828_, negedge _0560_)
    if (!_0560_) _3792_ <= 56'h000000204023d1;
    else _3792_ <= { _1989_[15:5], _1792_, _1989_[3:2], _1992_[8], _2168_[56:55], _2137_, _0297_, _0657_, _0698_, _1912_[29:15], _1592_, _1912_[13:10], _0188_, _1912_[8:2], _1915_[10:6] };
  assign { _2311_[55:48], _0863_, _2311_[46:16], _1623_, _2311_[14:0] } = _3792_;
  reg [1:0] _3793_;
  always_ff @(negedge _0241_, posedge _0467_)
    if (_0467_) _3793_ <= 2'h1;
    else _3793_ <= { _0298_, _0360_ };
  assign { _2312_[1], _0474_ } = _3793_;
  reg [5:0] _3794_;
  always_ff @(negedge _0134_, posedge _0690_)
    if (_0690_) _3794_ <= 6'h37;
    else _3794_ <= { _2170_[32:31], _1008_, _2170_[29:28], _1206_ };
  assign { _1014_, _1952_[141], _1621_, _1577_, _1320_, _1952_[137] } = _3794_;
  reg [58:0] _3795_;
  always_ff @(negedge _2026_[36], negedge _1139_)
    if (!_1139_) _3795_ <= 59'h7ffffffecd16719;
    else _3795_ <= { _2042_[11:1], _1336_, _2184_[13], _1630_, _2184_[11:6], _1740_, _2184_[4:0], _0907_, _0859_, _1135_, _1274_, _0741_, _0353_, _0249_, _0789_, _0801_, _0565_, _1993_[9:6], _1041_, _1993_[4:0], _0576_, _0844_, _1713_, _1822_, _0335_, _1834_, _2186_[3:2], _0932_, _0694_, _0666_, _0766_, _0046_ };
  assign { _1951_[116:105], _1560_, _1951_[103:88], _1910_[9:3], _1951_[80:58] } = _3795_;
  reg [30:0] _3796_;
  always_ff @(negedge _2118_[95], posedge _1133_)
    if (_1133_) _3796_ <= 31'h086d4a90;
    else _3796_ <= { _2004_[10:6], _1387_, _2018_[58:56], _0397_, _1640_, _0394_, _0763_, _0379_, _0573_, _0158_, _0949_, _1491_, _0047_, _0848_, _0005_, _0901_, _0296_, _1834_, _0149_, _0249_, _0758_, _1368_, _1627_, _0287_, _0144_ };
  assign { _2313_[30:22], _1782_, _2313_[20:0] } = _3796_;
  reg [29:0] _3797_;
  always_ff @(posedge _2050_[8], posedge _1148_)
    if (_1148_) _3797_ <= 30'h2ee0f5d2;
    else _3797_ <= { _0925_, _1939_[12:8], _0501_, _1939_[6], _1306_, _2000_[4], _1478_, _0042_, _0185_, _0338_, _0071_, _0913_, _1424_, _0772_, _0531_, _2003_[10:9], _1126_, _1631_, _2003_[6:3], _1372_, _1217_, _2003_[0] };
  assign { _2314_[29:22], _1946_[13:9], _2314_[16:6], _2239_, _2314_[4:0] } = _3797_;
  reg [133:0] _3798_;
  always_ff @(negedge _1165_, negedge _1656_)
    if (!_1656_) _3798_ <= 134'h0000000000000000000000000000000000;
    else _3798_ <= { _1952_[182:180], _0422_, _2058_[95:92], _1288_, _2058_[90:60], _1427_, _2058_[58:0], _1971_[25:19], _0922_, _1971_[17:13], _1525_, _1971_[11:0], _0325_, _0221_, _2312_[1], _0474_, _1966_[4], _0818_, _1966_[2], _0522_ };
  assign { _2315_[133:73], _1584_, _2315_[71:28], _2247_, _2315_[26:0] } = _3798_;
  reg [40:0] _3799_;
  always_ff @(negedge _0127_, negedge _0356_)
    if (!_0356_) _3799_ <= 41'h1ffc3f35d63;
    else _3799_ <= { _2112_[36:28], _1666_, _2112_[26:15], _0262_, _2112_[13:12], _1604_, _2112_[10:6], _0410_, _2112_[4:0], _0189_, _0127_, _0356_, _0101_ };
  assign { _2262_[56:54], _1690_, _2262_[52], _2025_[43:40], _1785_, _2025_[38:34], _1510_, _2025_[32:27], _0896_, _2025_[25], _1556_, _0114_, _0319_, _2041_[32:31], _1755_, _2041_[29:24], _0233_, _0499_, _2114_[25:23] } = _3799_;
  reg [6:0] _3800_;
  always_ff @(posedge _0287_, negedge _2047_[45])
    if (!_2047_[45]) _3800_ <= 7'h57;
    else _3800_ <= _2029_[38:32];
  assign { _2316_[6], _1582_, _2316_[4:2], _1605_, _2316_[0] } = _3800_;
  always_ff @(posedge _0585_, posedge _1514_)
    if (_1514_) _0479_ <= 1'h0;
    else _0479_ <= _1967_[12];
  reg [46:0] _3802_;
  always_ff @(posedge _0347_, negedge _1634_)
    if (!_1634_) _3802_ <= 47'h0000620a8675;
    else _3802_ <= { _2295_[22:12], _0750_, _2295_[10:4], _0057_, _1121_, _1862_, _1418_, _1228_, _0215_, _2155_[11:2], _1871_, _2155_[0], _0221_, _1481_, _0149_, _2133_[6:1], _1727_ };
  assign { _2317_[46:43], _2250_[70:42], _1749_, _2250_[40:33], _2317_[4:0] } = _3802_;
  reg [18:0] _3803_;
  always_ff @(posedge _1838_, negedge _2001_[104])
    if (!_2001_[104]) _3803_ <= 19'h2264f;
    else _3803_ <= { _2053_[36:28], _1667_, _2053_[26:21], _1211_, _0752_, _0134_ };
  assign { _2236_[22:19], _2215_[7:2], _1559_, _2213_[23:18], _2236_[5:4] } = _3803_;
  reg [6:0] _3804_;
  always_ff @(negedge _0435_, negedge _0041_)
    if (!_0041_) _3804_ <= 7'h45;
    else _3804_ <= { _2316_[6], _1582_, _2316_[4:2], _0510_, _0447_ };
  assign _2229_[37:31] = _3804_;
  reg [18:0] _3805_;
  always_ff @(posedge _2006_[3], negedge _1132_)
    if (!_1132_) _3805_ <= 19'h31bdb;
    else _3805_ <= { _1942_[16:15], _1279_, _1942_[13:10], _1619_, _1942_[8:7], _1602_, _0031_, _1077_, _0248_, _1684_, _2028_[3], _1326_, _2028_[1], _0598_ };
  assign { _0494_, _1930_[17:0] } = _3805_;
  reg [8:0] _3806_;
  always_ff @(posedge _0043_, posedge _1075_)
    if (_1075_) _3806_ <= 9'h076;
    else _3806_ <= { _2139_[35:32], _1354_, _1054_, _2139_[29:27] };
  assign _1956_[10:2] = _3806_;
  reg [12:0] _3807_;
  always_ff @(posedge _0811_, posedge _2157_[16])
    if (_2157_[16]) _3807_ <= 13'h0610;
    else _3807_ <= { _2093_[87:77], _1591_, _2093_[75] };
  assign { _1900_[62:59], _0498_, _1900_[57:54], _0066_, _1900_[52:50] } = _3807_;
  reg [14:0] _3808_;
  always_ff @(posedge _0354_, negedge _1098_)
    if (!_1098_) _3808_ <= 15'h2273;
    else _3808_ <= { _0811_, _1729_, _0064_, _1638_, _0369_, _0273_, _0302_, _0489_, _0488_, _0820_, _1845_, _0454_, _0445_, _0844_, _1713_ };
  assign { _2318_[14:7], _2253_[6:5], _2318_[4], _1877_, _2318_[2:0] } = _3808_;
  reg [49:0] _3809_;
  always_ff @(negedge _0463_, negedge _0690_)
    if (!_0690_) _3809_ <= 50'h3ffffe3eb97a2;
    else _3809_ <= { _1893_[10:7], _1034_, _1893_[5], _1070_, _2245_[79], _1313_, _0624_, _2141_[22:19], _2245_[72:70], _1984_[46:39], _1714_, _1984_[37:36], _0251_, _1984_[34:15], _2245_[37] };
  assign { _1979_[56:55], _1658_, _1979_[53], _1268_, _1979_[51:43], _1002_, _1979_[41:22], _0790_, _1979_[20:16], _1562_, _1979_[14:9], _1616_, _1979_[7] } = _3809_;
  reg [10:0] _3810_;
  always_ff @(posedge _2025_[40], posedge _0775_)
    if (_0775_) _3810_ <= 11'h1b9;
    else _3810_ <= { _2091_[11], _2014_[17:15], _1014_, _1952_[141], _1621_, _1577_, _1320_, _1952_[137], _0189_ };
  assign { _1964_[52], _1795_, _1964_[50:48], _1016_, _1964_[46:45], _0492_, _1964_[43], _1706_ } = _3810_;
  reg [167:0] _3811_;
  always_ff @(posedge _2066_[8], posedge _2318_[11])
    if (_2318_[11]) _3811_ <= 168'h000000000000000000000000000000000000000000;
    else _3811_ <= { _2148_[15:12], _0027_, _0560_, _0683_, _2125_[48:44], _0845_, _2125_[42:13], _1277_, _2125_[11:0], _0290_, _2133_[6:1], _1727_, _0202_, _0429_, _0683_, _0367_, _0718_, _1558_, _2219_[9:8], _0657_, _2171_, _0997_, _0814_, _0359_, _1046_, _2157_, _0979_, _0763_, _0208_, _0665_, _0712_, _2269_[12], _0892_, _2269_[10:8], _1050_, _0329_, _1813_, _2269_[4:0], _1457_, _1399_, _1711_, _1035_, _1967_[21:15], _1668_, _1967_[13:10], _1321_, _0473_, _1967_[7:0], _0306_, _0340_, _0731_, _0537_, _1112_ };
  assign { _2319_[167:35], _2243_[12:9], _2319_[30:0] } = _3811_;
  reg [4:0] _3812_;
  always_ff @(posedge _0287_, posedge _0907_)
    if (_0907_) _3812_ <= 5'h1a;
    else _3812_ <= { _1488_, _2040_[6:3] };
  assign _1992_[4:0] = _3812_;
  reg [14:0] _3813_;
  always_ff @(posedge _0361_, posedge _0594_)
    if (_0594_) _3813_ <= 15'h5543;
    else _3813_ <= { _2291_[14:11], _1628_, _2291_[9:2], _0259_, _0317_ };
  assign { _2320_[14:12], _0583_, _2320_[10:0] } = _3813_;
  reg [52:0] _3814_;
  always_ff @(posedge _0116_, posedge _0111_)
    if (_0111_) _3814_ <= 53'h0000005f1aab78;
    else _3814_ <= { _1984_[39], _1714_, _1984_[37:36], _0251_, _1984_[34:15], _0379_, _2000_[20:19], _0564_, _2000_[17:14], _0925_, _1939_[12:8], _0501_, _1939_[6], _1306_, _2000_[4:3], _1632_, _1373_, _2000_[0], _0125_, _1786_, _0402_, _1397_, _1569_, _1970_[5] };
  assign { _2321_[52], _1909_[39:35], _0254_, _1909_[33:25], _2204_[2], _1672_, _2321_[34:17], _1848_, _2321_[15], _1789_, _2321_[13:1], _2277_ } = _3814_;
  reg [12:0] _3815_;
  always_ff @(negedge _2047_[2], posedge _0033_)
    if (_0033_) _3815_ <= 13'h0619;
    else _3815_ <= { _2203_[10], _1571_, _2203_[8], _1938_[8:5], _0131_, _2203_[2], _0788_, _0479_, _0218_, _0490_ };
  assign _1955_[13:1] = _3815_;
  reg [68:0] _3816_;
  always_ff @(posedge _0274_, posedge _0731_)
    if (_0731_) _3816_ <= 69'h000000000000000000;
    else _3816_ <= { _2192_[32:24], _0298_, _0267_, _1639_, _1555_, _0287_, _0677_, _0843_, _0627_, _0020_, _0993_, _0403_, _0333_, _1486_, _0944_, _0071_, _0548_, _2015_[20:2], _1369_, _2015_[0], _0505_, _1116_, _0609_, _0134_, _1784_, _1956_[18:15], _0506_, _1956_[13:12], _0671_, _2117_[8:6], _0432_, _2117_[4:1], _2213_[3], _0802_ };
  assign { _2322_[68:57], _0073_, _2322_[55:38], _2249_[40:27], _1652_, _1241_, _2249_[24:7], _2322_[3:0] } = _3816_;
  reg [33:0] _3817_;
  always_ff @(negedge _0481_, negedge _1955_[18])
    if (!_1955_[18]) _3817_ <= 34'h030f7eb6b;
    else _3817_ <= { _2224_[14:1], _1172_, _0352_, _0357_, _0773_, _2135_, _0804_, _0241_, _1077_, _0248_, _1684_, _2028_[3], _1326_, _2028_[1] };
  assign { _1948_, _2323_[23:16], _1297_, _2323_[14:0] } = _3817_;
  reg [42:0] _3818_;
  always_ff @(posedge _0022_, negedge _0586_)
    if (!_0586_) _3818_ <= 43'h7fff4886388;
    else _3818_ <= { _1951_[157:151], _1276_, _1951_[149:144], _1042_, _1951_[142:139], _0356_, _0857_, _0531_, _0238_, _0633_, _0162_, _1959_[7], _1202_, _0226_, _0194_, _1964_[67], _0364_, _1888_[13], _0036_, _0706_, _1888_[10:5], _0673_, _1964_[55], _1679_ };
  assign { _1994_[9:6], _0840_, _1994_[4:3], _0597_, _2048_[51:50], _1423_, _2048_[48:47], _2005_[10:8], _1327_, _2005_[6:4], _2048_[39:38], _1150_, _2048_[36], _1010_, _2048_[34:17] } = _3818_;
  always_ff @(negedge _0810_, posedge _1955_[3])
    if (_1955_[3]) _0935_ <= 1'h0;
    else _0935_ <= _0304_;
  reg [3:0] _3820_;
  always_ff @(posedge _0018_, negedge _0361_)
    if (!_0361_) _3820_ <= 4'h6;
    else _3820_ <= { _2199_[18:17], _0144_, _0065_ };
  assign { _1225_, _1141_, _0622_, _1986_[1] } = _3820_;
  reg [6:0] _3821_;
  always_ff @(posedge _1981_[11], posedge _0203_)
    if (_0203_) _3821_ <= 7'h7c;
    else _3821_ <= { _0334_, _1786_, _0402_, _1397_, _1569_, _1970_[5], _0128_ };
  assign { _1493_, _2020_[10:9], _0293_, _2020_[7:5] } = _3821_;
  reg [9:0] _3822_;
  always_ff @(negedge _0926_, posedge _0227_)
    if (_0227_) _3822_ <= 10'h123;
    else _3822_ <= { _2169_[50:45], _1793_, _2169_[43:41] };
  assign { _1900_[72:70], _0389_, _1900_[68:66], _0833_, _1305_, _1900_[63] } = _3822_;
  reg [5:0] _3823_;
  always_ff @(posedge _1677_, posedge _0573_)
    if (_0573_) _3823_ <= 6'h28;
    else _3823_ <= _2035_[11:6];
  assign { _1077_, _0248_, _1684_, _2028_[3], _1326_, _2028_[1] } = _3823_;
  reg [6:0] _3824_;
  always_ff @(negedge _0549_, posedge _1587_)
    if (_1587_) _3824_ <= 7'h63;
    else _3824_ <= { _1999_[107:105], _0228_, _0013_, _1865_, _1192_ };
  assign _1893_[44:38] = _3824_;
  assign _1886_[14] = _1620_;
  assign { _1887_[13], _1887_[9], _1887_[7] } = { _0852_, _1850_, _1537_ };
  assign { _1888_[12:11], _1888_[4:2], _1888_[0] } = { _0036_, _0706_, _0673_, _0059_, _0148_, _0479_ };
  assign { _1889_[12:11], _1889_[7:6] } = { _0596_, _1753_, _1624_, _1312_ };
  assign { _1890_[12], _1890_[10:9], _1890_[5:0] } = { _0588_, _0350_, _0716_, _1136_, _0238_, _0109_, _0306_, _0116_, _0238_ };
  assign _1891_[4:0] = { _0639_, _1009_, _0109_, _1283_, _0219_ };
  assign { _1893_[55:51], _1893_[48:45], _1893_[13:11], _1893_[6], _1893_[3:0] } = { _0766_, _0490_, _0526_, _1609_, _0241_, _0771_, _0807_, _0894_, _0551_, _0702_, _1402_, _1153_, _1034_, _1374_, _1787_, _0126_, _1328_ };
  assign { _1894_[47:46], _1894_[40], _1894_[37:19], _1894_[2:0] } = { _0043_, _0213_, _0676_, _0445_, _0179_, _0496_, _0476_, _0054_, _0677_, _0349_, _1025_, _0298_, _1171_, _1218_, _0269_, _0476_, _0470_, _1733_, _1065_, _0390_, _1220_, _0886_, _0043_, _0944_, _0076_ };
  assign { _1895_[25], _1895_[19], _1895_[1:0] } = { _1111_, _1757_, _0281_, _1171_ };
  assign { _1896_[23], _1896_[11], _1896_[8], _1896_[5:0] } = { _1594_, _1712_, _0096_, _0030_, _0639_, _0359_, _0987_, _1626_, _1611_ };
  assign { _1897_[51], _1897_[26], _1897_[20] } = { _1665_, _1260_, _0037_ };
  assign { _1898_[53:39], _1898_[22], _1898_[16], _1898_[9] } = { _0405_, _0922_, _0062_, _1036_, _0381_, _0289_, _0636_, _0565_, _0398_, _1182_, _0884_, _0526_, _0599_, _1171_, _0858_, _1517_, _1593_, _0765_ };
  assign _1899_[2:0] = { _0079_, _0911_, _0303_ };
  assign { _1900_[78:77], _1900_[75], _1900_[73], _1900_[69], _1900_[65:64], _1900_[58], _1900_[53], _1900_[49:47], _1900_[36], _1900_[28:27], _1900_[25:22], _1900_[19:1] } = { _1760_, _0451_, _0191_, _1491_, _0389_, _0833_, _1305_, _0498_, _0066_, _0689_, _1409_, _1639_, _0767_, _0230_, _1833_, _1394_, _0384_, _0358_, _0334_, _0804_, _0080_, _0510_, _0596_, _1753_, _1889_[10:8], _1624_, _1312_, _1889_[5:0], _1018_, _0518_, _1820_ };
  assign { _1901_[73], _1901_[69:67], _1901_[62], _1901_[60], _1901_[58], _1901_[38:29], _1901_[27:18], _1901_[16], _1901_[13], _1901_[9], _1901_[4] } = { _0107_, _0465_, _0082_, _0092_, _1575_, _1370_, _1023_, _0225_, _1229_, _0133_, _1893_[44:38], _1623_, _0678_, _0198_, _1481_, _0827_, _0325_, _0271_, _1171_, _0548_, _0317_, _0555_, _0760_, _0879_, _1078_ };
  assign _1902_[28] = _1293_;
  assign { _1903_[35], _1903_[2:0] } = { _1213_, _1742_, _1555_, _1149_ };
  assign { _1904_[21:10], _1904_[1:0] } = { _1599_, _1893_[44:38], _0698_, _0821_, _1812_, _0971_, _0272_, _0001_ };
  assign _1905_[4] = _0077_;
  assign _1906_[0] = _0744_;
  assign { _1907_[24], _1907_[15], _1907_[13], _1907_[11], _1907_[9:8] } = { _1535_, _0900_, _1017_, _0011_, _0867_, _0134_ };
  assign { _1908_[37], _1908_[35], _1908_[20:17], _1908_[15], _1908_[12], _1908_[9], _1908_[6:0] } = { _1885_, _1270_, _0620_, _0875_, _0531_, _0117_, _0986_, _1564_, _0535_, _0016_, _1208_, _1491_, _0611_, _0421_, _1809_, _0652_ };
  assign { _1909_[34], _1909_[24:23], _1909_[21:20], _1909_[17:16], _1909_[14], _1909_[11:5], _1909_[1:0] } = { _0254_, _0539_, _0807_, _1290_, _1096_, _0237_, _0032_, _0561_, _1908_[39:38], _1885_, _1908_[36], _1270_, _1908_[34], _1048_, _1167_, _0607_ };
  assign _1910_[2:1] = { _0010_, _0304_ };
  assign { _1911_[7:5], _1911_[0] } = { _1284_, _0908_, _0573_, _1329_ };
  assign { _1912_[39:37], _1912_[35], _1912_[33], _1912_[31:30], _1912_[14], _1912_[9], _1912_[1] } = { _0289_, _0109_, _1019_, _1729_, _1564_, _0019_, _1183_, _1592_, _0188_, _0631_ };
  assign { _1913_[39:37], _1913_[30], _1913_[24:23], _1913_[9], _1913_[7:6], _1913_[4], _1913_[2:0] } = { _0134_, _0453_, _0442_, _1466_, _0567_, _1701_, _1821_, _1035_, _0642_, _0733_, _0234_, _1088_, _0454_ };
  assign { _1914_[39:33], _1914_[31:18], _1914_[16], _1914_[14:11], _1914_[9:1] } = { _0948_, _1868_, _1742_, _1827_, _0490_, _0204_, _0641_, _0440_, _0634_, _0848_, _0116_, _0411_, _0837_, _1629_, _1208_, _0419_, _0641_, _0232_, _0848_, _0872_, _1644_, _0096_, _1887_[14], _0852_, _1887_[12], _0477_, _1529_, _1348_, _0226_, _0598_, _1641_, out_data[1184], _0967_, _1641_, _0372_ };
  assign { _1915_[46:44], _1915_[12:11], _1915_[5:3], _1915_[1] } = { _0914_, _1725_, _0186_, _0103_, _1329_, _0452_, _0385_, _1165_, _0179_ };
  assign { _1916_[8], _1916_[5:3], _1916_[1:0] } = { _1139_, _1656_, _0873_, _0915_, _0631_, _1299_ };
  assign { _1917_[13:11], _1917_[9], _1917_[4], _1917_[2], _1917_[0] } = { _0287_, _0936_, _0642_, _1208_, _1731_, _1087_, _1363_ };
  assign { _1918_[10], _1918_[1] } = { _1295_, _0937_ };
  assign { _1919_[16], _1919_[6], _1919_[4:0] } = { _0557_, _1882_, _0904_, _1125_, _1025_, _0882_, _0856_ };
  assign { _1920_[21], _1920_[18], _1920_[15], _1920_[1:0] } = { _0056_, _1816_, _1168_, _1841_, _0299_ };
  assign _1923_[1:0] = { _1343_, _0342_ };
  assign _1924_[6:3] = { _0847_, _1630_, _0372_, _1380_ };
  assign { _1925_[6:5], _1925_[0] } = { _1138_, _0936_, _0134_ };
  assign { _1926_[4], _1926_[1] } = { _0614_, _1818_ };
  assign { _1927_[24:23], _1927_[21:20], _1927_[18], _1927_[5:3], _1927_[1:0] } = { _0069_, _0208_, _1046_, _0609_, _1565_, _0853_, _1343_, _1453_, _1447_, _0133_ };
  assign { _1928_[17], _1928_[11], _1928_[8:7], _1928_[5], _1928_[3:0] } = { _0244_, _0441_, _1170_, _0134_, _0592_, _0325_, _0014_, _0951_, _0565_ };
  assign { _1929_[27], _1929_[24:16], _1929_[14:5], _1929_[2:0] } = { _0355_, _0342_, _0071_, _0321_, _0700_, _0082_, _1360_, _1188_, _1589_, _0752_, _0873_, _0026_, _0315_, _0599_, _0480_, _0454_, _0315_, _0482_, _1761_, _1590_, _0046_, _0715_, _1486_ };
  assign { _1930_[27:23], _1930_[21:20], _1930_[18] } = { _1901_[56:53], _0228_, _0438_, _0297_, _0494_ };
  assign _1931_[1:0] = { _1720_, _0449_ };
  assign { _1932_[12:7], _1932_[5], _1932_[3], _1932_[1:0] } = { _1235_, _0269_, _1329_, _1607_, _1810_, _0123_, _0595_, out_data[416], _0430_, _0449_ };
  assign { _1933_[29], _1933_[17:16], _1933_[8], _1933_[5:4], _1933_[2:0] } = { out_data[544], _1258_, _0894_, _1244_, _0421_, _0152_, _1006_, _0846_, _0580_ };
  assign _1934_[3:0] = { _0335_, _0005_, _0882_, _0941_ };
  assign { _1935_[78], _1935_[71:67], _1935_[65:64], _1935_[61], _1935_[59:58], _1935_[55:48], _1935_[37:31], _1935_[29:27], _1935_[23:22], _1935_[20:19], _1935_[16], _1935_[14:0] } = { _1157_, _0044_, _1615_, _0342_, _0873_, _1657_, _0314_, _0599_, _0400_, _0103_, _0270_, _0873_, _0636_, _0563_, _0549_, _0146_, _0559_, _1484_, _1770_, _0546_, _1916_[6], _1656_, _0038_, _0198_, _0302_, _0490_, _0882_, _1424_, _1539_, _0206_, _0401_, _1478_, _1406_, _0558_, _0411_, _0338_, _0596_, _1753_, _1889_[10:8], _1624_, _1312_, _1889_[5:0] };
  assign { _1936_[54], _1936_[52:48], _1936_[43], _1936_[41], _1936_[39:10], _1936_[8:5], _1936_[3:0] } = { _1621_, _0348_, _1075_, _0940_, _1123_, _0651_, _1612_, _0418_, _1913_[36:31], _1466_, _1913_[29:25], _0567_, _1701_, _1913_[22:10], _1821_, _1913_[8], _0067_, _0103_, _1411_, _0191_, _0219_, _0801_, _1622_, _0488_, _0639_ };
  assign _1938_[4:1] = { _0609_, _0076_, _0241_, _0134_ };
  assign { _1939_[7], _1939_[5:4], _1939_[2:1] } = { _0501_, _1134_, _1225_, _0321_, _0116_ };
  assign { _1940_[37], _1940_[25], _1940_[23], _1940_[19:3], _1940_[1] } = { _1446_, _1696_, _1230_, _1901_[86:74], _0107_, _1901_[72:70], _0351_ };
  assign { _1941_[23:14], _1941_[0] } = { _1421_, _0489_, _0038_, _0115_, _0810_, _0338_, _1820_, _0043_, _1037_, _1567_, _0895_ };
  assign { _1942_[57:56], _1942_[53:48], _1942_[44], _1942_[38], _1942_[22:21], _1942_[19:17], _1942_[14], _1942_[9], _1942_[2:0] } = { _0111_, _0454_, _0004_, _0144_, _0317_, _0860_, _1362_, _0489_, _1285_, _1547_, _1512_, _0519_, _1139_, _0096_, _0279_, _1279_, _1619_, _0437_, _0562_, _0539_ };
  assign { _1943_[110], _1943_[88:83], _1943_[74], _1943_[67], _1943_[63], _1943_[44:38], _1943_[24], _1943_[4], _1943_[0] } = { _1768_, _0047_, _0678_, _0183_, _0094_, _0619_, _0253_, _1082_, _1504_, _1724_, _0287_, _1720_, _0105_, _1228_, _0585_, _0306_, _1453_, _1498_, _0647_, _0991_ };
  assign { _1944_[34:30], _1944_[4:1] } = { _0893_, _1270_, _0259_, _1453_, _0904_, _0799_, _0206_, _1876_, _0143_ };
  assign { _1945_[4:3], _1945_[1] } = { _0631_, _1077_, _0442_ };
  assign _1946_[0] = _1462_;
  assign { _1947_[13:12], _1947_[5], _1947_[2:0] } = { _0764_, _0206_, _1267_, _1646_, _0522_, _0149_ };
  assign _1949_[4:0] = { _1883_, _0366_, _0372_, _0982_, _0025_ };
  assign _1950_[195:164] = out_data[1311:1280];
  assign { _1951_[215:170], _1951_[158], _1951_[150], _1951_[143], _1951_[138:137], _1951_[133:131], _1951_[127:124], _1951_[122], _1951_[118:117], _1951_[104], _1951_[87:81], _1951_[57:34], _1951_[32], _1951_[30], _1951_[5], _1951_[1:0] } = { _1897_[47:27], _1260_, _1897_[25:21], _0037_, _1897_[19:4], _0228_, _0625_, _1255_, _1276_, _1042_, _0124_, _0929_, _0505_, _0423_, _0087_, _0235_, _0917_, _0917_, out_data[544], _1122_, _1609_, _0080_, _1560_, _1910_[9:3], _0285_, _0868_, _0977_, _1429_, _0413_, _0879_, _1486_, _0334_, _0032_, _0412_, _0118_, _1085_, _0529_, _0217_, _1880_, _0442_, _0325_, _1178_, _0015_, _1561_, _0964_, _1831_, _1555_, _1606_, _1412_, _1496_, _0382_, _0800_, _1371_ };
  assign { _1952_[213], _1952_[205], _1952_[183], _1952_[176], _1952_[164], _1952_[156:142], _1952_[140:138], _1952_[136:60], _1952_[44:43], _1952_[41], _1952_[16], _1952_[11], _1952_[6], _1952_[3:0] } = { _1083_, _1246_, _1389_, _0344_, _1194_, _0228_, _1758_, _1659_, _0292_, _0054_, _1144_, _1777_, _0420_, _0357_, _0145_, _0044_, _0701_, _1021_, _0804_, _1014_, _1621_, _1577_, _1320_, _1648_, _0278_, _0811_, _0855_, _1657_, _0028_, _1780_, _0683_, _1362_, _0175_, _1301_, _0029_, _1433_, _1177_, _1138_, _0797_, _1892_, _0939_, _0362_, _0324_, _0379_, _1215_, _1232_, _1494_, _0803_, _1586_, _1385_, _1118_, out_data[1888], _1554_, _0217_, _1044_ };
  assign { _1953_[28:25], _1953_[7], _1953_[5:0] } = { _1935_[75:72], _1428_, _0611_, _1463_, _0835_, _1033_, _1599_, _1664_ };
  assign { _1954_[11], _1954_[8] } = { _1872_, out_data[1952] };
  assign { _1955_[30:26], _1955_[19], _1955_[17], _1955_[15], _1955_[0] } = { _1952_[52:48], _0072_, _1853_, _1487_, _0217_ };
  assign { _1956_[23], _1956_[21:19], _1956_[14], _1956_[11], _1956_[1:0] } = { _1618_, _1642_, _1629_, _0017_, _0506_, _0828_, _0218_, _0273_ };
  assign _1957_[13:2] = { _1904_[36:31], _0950_, _1190_, _0933_, _0358_, _0102_, _1870_ };
  assign _1958_[3:0] = { _0661_, _0875_, _0359_, _1137_ };
  assign { _1959_[9:8], _1959_[6:5], _1959_[2:0] } = { _0633_, _0162_, _1202_, _1431_, _1145_, _1089_, _0948_ };
  assign _1960_[34:3] = out_data[639:608];
  assign _1961_[0] = _0000_;
  assign { _1962_[34:12], _1962_[4], _1962_[0] } = { out_data[1276:1254], _1261_, _0228_ };
  assign _1963_[59:28] = out_data[511:480];
  assign { _1964_[76], _1964_[73], _1964_[66:56], _1964_[54:53], _1964_[51], _1964_[47], _1964_[44], _1964_[42:33], _1964_[30], _1964_[26:22], _1964_[6:0] } = { _1452_, _1647_, _0364_, _1888_[13], _0036_, _0706_, _1888_[10:5], _0673_, _1679_, _1617_, _1795_, _1016_, _0492_, _1706_, _0890_, _1084_, _1831_, _0843_, _0721_, _0960_, _0480_, _0268_, _1381_, _1156_, _1264_, _1299_, _0568_, _0915_, _0355_, _1092_, _0232_, _0615_, out_data[864], _0934_, _0018_, _1394_ };
  assign _1965_[77:46] = out_data[319:288];
  assign { _1966_[64:45], _1966_[41:40], _1966_[33], _1966_[26:25], _1966_[18], _1966_[13:10], _1966_[8:5], _1966_[3], _1966_[1:0] } = { _1052_, _0447_, _0096_, _1275_, _1299_, _0062_, _1207_, _1580_, _1876_, _0189_, _0068_, _1043_, _1933_[13:9], _1244_, _1933_[7:6], _1236_, _1174_, _0990_, _0988_, _1879_, _0528_, _0540_, _1864_, _1186_, _1505_, _0631_, _1744_, _0259_, _1549_, _0818_, _0807_, _0636_ };
  assign { _1967_[77:36], _1967_[22], _1967_[14], _1967_[9:8] } = { _1920_[16], _1168_, _1920_[14], _0241_, _0752_, _1079_, _0756_, _0082_, _0586_, _1063_, _0025_, _1913_[36:31], _1466_, _1913_[29:25], _0567_, _1701_, _1913_[22:10], _1821_, _1913_[8], _1259_, _0301_, _1123_, _1668_, _1321_, _0473_ };
  assign { _1968_[51], _1968_[49], _1968_[13] } = { _0719_, _1022_, _0142_ };
  assign { _1969_[35], _1969_[28], _1969_[7:0] } = { _0677_, _0985_, _0453_, _1266_, _0096_, _0529_, _0752_, _1283_, _0625_, _0065_ };
  assign { _1970_[19], _1970_[15:14], _1970_[10:6], _1970_[4:0] } = { _1253_, _1210_, _1682_, _0159_, _1786_, _0402_, _1397_, _1569_, _0716_, _0907_, _0206_, _0241_, _0071_ };
  assign { _1971_[18], _1971_[12] } = { _0922_, _1525_ };
  assign { _1972_[21], _1972_[10:0] } = { _1687_, _1310_, _0636_, _0678_, _0993_, _0403_, _0589_, _0739_, _0918_, _0101_, _0639_, _0518_ };
  assign { _1973_[23:21], _1973_[18:0] } = { _0504_, _1597_, _0684_, _1970_[51:39], _0464_, _1235_, _1374_, _0356_, _0999_, _0194_ };
  assign _1974_[1] = _0155_;
  assign { _1975_[53], _1975_[51:23] } = { _1790_, _1926_[30:5], _0614_, _1926_[3:2] };
  assign { _1976_[74:71], _1976_[57], _1976_[33], _1976_[25], _1976_[22:20], _1976_[15], _1976_[13:11], _1976_[8], _1976_[6], _1976_[4] } = { _0189_, _0033_, _0065_, _0018_, _1797_, _0100_, _1341_, _0121_, _0563_, _0591_, _1335_, _0172_, _0120_, _1568_, _0604_, _0945_, _0602_ };
  assign { _1977_[74:26], _1977_[23:0] } = { _1889_[2], _1976_[70:58], _1797_, _1976_[56:34], _0100_, _1976_[32:26], _1341_, _1976_[24:23], _1243_, _1384_, _1669_, _0256_, _0116_, _1203_, _0983_, _1046_, _0915_, _0019_, _0227_, _0356_, _1621_, _0155_, _1974_[0], _1527_, _1374_, _0217_, _0043_, _0134_, _0069_, _0311_, _0134_, _0046_ };
  assign _1978_[48:14] = { _1446_, _1940_[36:26], _1696_, _1940_[24], _1230_, _1940_[22:20], _1901_[86:74], _0107_, _1901_[72:70] };
  assign { _1979_[58:57], _1979_[54], _1979_[52], _1979_[42], _1979_[21], _1979_[15], _1979_[8], _1979_[6:0] } = { _1976_[37:36], _1658_, _1268_, _1002_, _0790_, _1562_, _1616_, _1621_, _0238_, _0071_, _0401_, _0287_, _0857_, _0049_ };
  assign { _1980_[5], _1980_[3] } = { _1367_, _1681_ };
  assign { _1981_[23:12], _1981_[8:7], _1981_[1:0] } = { _0025_, _0238_, _0617_, _0625_, _0025_, _0151_, _0043_, _0469_, _1951_[33], _1412_, _1951_[31], _1496_, _0299_, _0223_, _1794_, _0194_ };
  assign { _1982_[23:22], _1982_[15], _1982_[5:0] } = { _1381_, _1520_, _1534_, _1287_, _0174_, _0343_, _0383_, _0265_, _0453_ };
  assign _1983_[25:10] = { _1928_[24:18], _0244_, _1928_[16:12], _0441_, _1928_[10:9] };
  assign { _1984_[38], _1984_[35], _1984_[14:0] } = { _1714_, _0251_, _0243_, _0739_, _1153_, _1893_[10:7], _1034_, _1893_[5:4], _1374_, _1787_, _0126_, _1328_, _0254_ };
  assign _1985_[1] = _1692_;
  assign { _1986_[11:2], _1986_[0] } = { _0350_, _0716_, _0565_, _0572_, _1374_, _1527_, _0518_, _1225_, _1141_, _0622_, _0068_ };
  assign { _1987_[51], _1987_[47], _1987_[30], _1987_[22] } = { _1596_, _1839_, _0693_, _0798_ };
  assign { _1988_[50], _1988_[48], _1988_[45], _1988_[42], _1988_[37], _1988_[35], _1988_[26:25], _1988_[23], _1988_[21], _1988_[18:0] } = { _0291_, _1383_, _1697_, _0277_, _0130_, _0725_, _1406_, _1175_, _0921_, _1819_, _0102_, _0697_, _0690_, _1964_[67], _0364_, _1888_[13], _0036_, _0706_, _1888_[10:5], _0673_, _1964_[55], _1679_, _0589_, _0096_ };
  assign { _1989_[32], _1989_[4], _1989_[1:0] } = { _1344_, _1792_, _0134_, _0311_ };
  assign { _1990_[54], _1990_[52], _1990_[44], _1990_[22], _1990_[15], _1990_[12] } = { _1811_, _1413_, _1764_, _1074_, _0928_, _0495_ };
  assign { _1991_[46:45], _1991_[42:0] } = { _1193_, _1553_, _0219_, _0887_, _0359_, _0642_, _0019_, _1951_[169:159], _1255_, _1951_[157:151], _1276_, _1951_[149:144], _1042_, _1951_[142:139], _0124_, _0929_, _1951_[136:134], _0678_, _1007_ };
  assign { _1992_[55:9], _1992_[7:5] } = { _1989_[48:33], _1344_, _1989_[31:5], _1792_, _1989_[3:2], _0189_, _0221_, _0566_ };
  assign _1993_[5] = _1041_;
  assign { _1994_[5], _1994_[2:0] } = { _0840_, _0597_, _0594_, _0999_ };
  assign { _1995_[13], _1995_[5], _1995_[0] } = { _0224_, _1242_, _1011_ };
  assign { _1996_[17:5], _1996_[3:0] } = { in_data[836:826], _1203_, _1716_, _1365_, _0104_, _1476_, _1467_ };
  assign _1998_[29] = _1325_;
  assign { _1999_[119], _1999_[99], _1999_[75], _1999_[66], _1999_[31] } = { _1109_, _1030_, _1817_, _0574_, _1303_ };
  assign { _2000_[139:124], _2000_[107], _2000_[99], _2000_[97], _2000_[91], _2000_[85], _2000_[79:60], _2000_[49], _2000_[45:43], _2000_[34], _2000_[30], _2000_[26:21], _2000_[18], _2000_[13:5], _2000_[2:1] } = { _1908_[10], _0535_, _1908_[8:7], _0363_, _0325_, _0210_, _0155_, _1974_[0], _0566_, _1007_, _0096_, _1951_[33], _1412_, _1951_[31], _1496_, _1361_, _1506_, _0113_, _0313_, _0737_, _0401_, _0105_, _0082_, _0152_, _0642_, _0108_, _0572_, _0317_, _0057_, _1951_[33], _1412_, _1951_[31], _1496_, _1225_, _1141_, _0622_, _1986_[1], _0095_, _1393_, _0241_, _1570_, _1314_, _1419_, _0391_, _1747_, _1307_, _1318_, _0097_, _1009_, _0502_, _0401_, _0125_, _0564_, _0925_, _1939_[12:8], _0501_, _1939_[6], _1306_, _1632_, _1373_ };
  assign { _2001_[137], _2001_[112], _2001_[110], _2001_[108:107], _2001_[102], _2001_[98], _2001_[96], _2001_[85], _2001_[72], _2001_[70:0] } = { _0211_, _0752_, _1323_, _1309_, _1081_, _1351_, _1353_, _1359_, _0998_, _1765_, _0719_, _1968_[50], _1022_, _1968_[48:14], _0142_, _1968_[12:0], _0287_, _0290_, _0015_, _0368_, _0278_, _0434_, _1985_[11:2], _1692_, _1985_[0], _0521_ };
  assign { _2002_[31:28], _2002_[25:7] } = { _1677_, _0409_, _1804_, _1386_, _1381_, _1520_, _1982_[21:16], _1534_, _1982_[14:6], _1287_ };
  assign { _2003_[8:7], _2003_[2:1] } = { _1126_, _1631_, _1372_, _1217_ };
  assign _2004_[5:0] = { _1387_, _0581_, _0572_, _0318_, _0359_, _0117_ };
  assign { _2005_[7], _2005_[3:0] } = { _1327_, _0189_, _0320_, _0278_, _0988_ };
  assign { _2006_[8:7], _2006_[5], _2006_[2:0] } = { _1254_, _0468_, _0404_, _1931_[3], _1308_, _0513_ };
  assign _2007_[0] = _0103_;
  assign _2008_[2:1] = { _1531_, _1068_ };
  assign { _2009_[3], _2009_[1:0] } = { _1805_, _0819_, _1807_ };
  assign _2010_[0] = _0240_;
  assign { _2011_[27], _2011_[5] } = { _1044_, _0181_ };
  assign { _2012_[27], _2012_[21:20], _2012_[1:0] } = { _1625_, _1678_, _1222_, _1613_, _0082_ };
  assign { _2013_[9], _2013_[6:5] } = { _1857_, _1829_, _1040_ };
  assign _2014_[9:0] = { _1988_[54:51], _0291_, _1988_[49], _1383_, _1988_[47:46], _0097_ };
  assign { _2015_[21], _2015_[1] } = { _0548_, _1369_ };
  assign _2016_[5:0] = { _0145_, _0122_, _0042_, _1449_, _0594_, _0781_ };
  assign { _2017_[60], _2017_[36], _2017_[32], _2017_[13] } = { _1364_, _1410_, _0414_, _1442_ };
  assign { _2018_[65:59], _2018_[55:54], _2018_[52:0] } = { _0920_, _2004_[10:6], _1387_, _0397_, _1640_, _0023_, _1449_, _0191_, _1265_, _0589_, _0907_, _0620_, _0206_, _0311_, _2000_[20:19], _0564_, _2000_[17:14], _0925_, _1939_[12:8], _0501_, _1939_[6], _1306_, _2000_[4:3], _1632_, _1373_, _2000_[0], _0795_, _0108_, _1203_, _0854_, _0986_, _1908_[14:13], _1564_, _1908_[11:10], _0535_, _1908_[8:7], _0984_, _0477_, _1329_, _0716_, _0600_, _0146_, _0572_, _0856_, _0134_, _0692_ };
  assign { _2019_[65:59], _2019_[56], _2019_[36:6], _2019_[4:0] } = { _1970_[42:38], _0117_, _0272_, _1636_, _0070_, _1920_[31:22], _0056_, _1920_[20:19], _1816_, _1920_[17:16], _1168_, _1920_[14:2], _1655_, _0452_, _0095_, _0318_, _0873_ };
  assign { _2020_[27:11], _2020_[8], _2020_[4:0] } = { _1985_[5:2], _1692_, _0235_, _0275_, _0316_, _0272_, _0325_, _1046_, _0324_, _1322_, _0254_, _0469_, _0044_, _1493_, _0293_, _0044_, _0608_, _0178_, _0726_, _0715_ };
  assign { _2021_[17], _2021_[12] } = { _0688_, _1189_ };
  assign { _2022_[21:9], _2022_[5], _2022_[2] } = { _0208_, _0235_, _0986_, _1908_[14:13], _1564_, _1908_[11:10], _0535_, _1908_[8:7], _1561_, _0619_, _1160_, _1069_ };
  assign { _2023_[11:10], _2023_[6] } = { _1469_, _1408_, _0327_ };
  assign { _2024_[11], _2024_[1:0] } = { _1825_, _0274_, _0016_ };
  assign { _2025_[39], _2025_[33], _2025_[26], _2025_[24:0] } = { _1785_, _1510_, _0896_, _0290_, _0133_, _0627_, _0043_, _0656_, _0716_, _0145_, _0752_, _1993_[9:6], _1041_, _1993_[4:0], _0627_, _0057_, _0383_, _0620_, _0281_, _0259_, _0058_ };
  assign { _2026_[33], _2026_[10], _2026_[6:0] } = { _0842_, _1097_, _0116_, _0097_, _1621_, _0111_, _0221_, _0176_, _0309_ };
  assign { _2027_[8], _2027_[4], _2027_[0] } = { _0889_, _0260_, _1107_ };
  assign { _2028_[10:4], _2028_[2], _2028_[0] } = { _2000_[123:122], _0690_, _1283_, _1077_, _0248_, _1684_, _1326_, _0489_ };
  assign { _2029_[43], _2029_[29], _2029_[18], _2029_[16], _2029_[10] } = { _1801_, _1012_, _1357_, _1440_, _1115_ };
  assign { _2030_[45], _2030_[41], _2030_[15] } = { _0705_, _1598_, _1685_ };
  assign { _2031_[65], _2031_[63:62], _2031_[54], _2031_[52], _2031_[50], _2031_[46:34], _2031_[30], _2031_[22], _2031_[18], _2031_[16:15], _2031_[2:0] } = { _0328_, _0007_, _1699_, _1806_, _0206_, _1800_, _1991_[55:47], _1193_, _1553_, _1991_[44:43], _1788_, _0514_, _1887_[16], _1101_, _1814_, _1509_, _0401_, _0235_ };
  assign { _2032_[53:32], _2032_[25], _2032_[12], _2032_[9], _2032_[0] } = { _1527_, _0228_, _0149_, _1265_, _0272_, _0915_, _2008_[14:3], _1531_, _1068_, _2008_[0], _1028_, _1826_, _0606_, _1754_, _0617_ };
  assign { _2033_[21], _2033_[5] } = { _1783_, _1407_ };
  assign _2034_[14:0] = { _0000_, _0700_, _0153_, _0634_, _0739_, _0185_, _0146_, _0304_, _0278_, _0238_, _0697_, _0196_, _0589_, _0572_, _0529_ };
  assign { _2035_[18:17], _2035_[15], _2035_[1:0] } = { _1455_, _1507_, _1674_, _0320_, _0795_ };
  assign { _2036_[13:12], _2036_[2] } = { _0509_, _0236_, _1715_ };
  assign { _2037_[25], _2037_[20] } = { _1823_, _1515_ };
  assign { _2038_[47], _2038_[45], _2038_[42:41], _2038_[24], _2038_[10:2] } = { _1039_, _0092_, _0630_, _0407_, _1060_, _2034_[23:15] };
  assign _2039_[10:0] = { _1417_, _0566_, _1464_, _0581_, _0455_, _0042_, _0518_, _0241_, _1368_, _0795_, _1550_ };
  assign { _2040_[35:21], _2040_[10:9], _2040_[7], _2040_[2:0] } = { in_data[1342:1333], _0043_, _0275_, _0043_, _0082_, _0317_, _0618_, _1485_, _1488_, _0096_, _0690_, _0068_ };
  assign { _2041_[35:33], _2041_[30], _2041_[23:0] } = { _1556_, _0114_, _0319_, _1755_, _0733_, _0915_, _0316_, _0189_, _0194_, _2001_[111], _1323_, _2001_[109], _1309_, _1081_, _2001_[106:103], _1351_, _2001_[101:99], _1353_, _2001_[97], _1359_, _0152_, _1000_, _0356_ };
  assign _2042_[0] = _1532_;
  assign _2043_[1:0] = { _0605_, _1009_ };
  assign { _2044_[5], _2044_[0] } = { _0668_, _1461_ };
  assign _2045_[4:0] = { _2012_[43:40], _0524_ };
  assign { _2046_[21:7], _2046_[5], _2046_[3] } = { _2038_[27:25], _1060_, _2038_[23:21], _0116_, _0354_, _0522_, _0187_, _0249_, _0217_, _0242_, _0193_, _1756_, _1094_ };
  assign { _2047_[79], _2047_[57], _2047_[13], _2047_[4], _2047_[1] } = { _1445_, _0850_, _1617_, _0679_, _0954_ };
  assign { _2048_[83:52], _2048_[49], _2048_[46:40], _2048_[37], _2048_[35], _2048_[16:0] } = { _1969_[34:29], _0985_, _1969_[27:15], _0383_, _0186_, _1127_, _0133_, _1994_[9:6], _0840_, _1994_[4:3], _0597_, _1423_, _2005_[10:8], _1327_, _2005_[6:4], _1150_, _1010_, _0192_, _2023_[13:12], _1469_, _1408_, _2023_[9:7], _0327_, _2023_[5:0], _0425_, _0091_ };
  assign { _2049_[71], _2049_[68:0] } = { _1121_, _2030_[66:46], _0705_, _2030_[44:42], _1598_, _2030_[40:16], _1685_, _2030_[14:0], _0995_, _0082_ };
  assign { _2050_[4], _2050_[1] } = { _1164_, _1296_ };
  assign _2051_[8:0] = { _1056_, _0121_, _0043_, _0642_, _0161_, _1360_, _0135_, _0146_, _0144_ };
  assign { _2052_[30:29], _2052_[16] } = { _0252_, _0331_, _0777_ };
  assign { _2053_[27], _2053_[20], _2053_[14], _2053_[10:0] } = { _1667_, _1695_, _1185_, _0129_, _0141_, _0152_, _0254_, _1044_, _1066_, _0116_, _0058_, _0071_, _0161_, _0340_ };
  assign { _2054_[38:35], _2054_[30], _2054_[18], _2054_[15], _2054_[8], _2054_[1:0] } = { _2039_[13:11], _1417_, _1683_, _1538_, _1029_, _1337_, _1633_, _0156_ };
  assign _2055_[3] = _1415_;
  assign _2056_[0] = _0510_;
  assign _2057_[0] = _1023_;
  assign { _2058_[91], _2058_[59] } = { _1288_, _1427_ };
  assign { _2059_[88], _2059_[75], _2059_[70], _2059_[66], _2059_[54], _2059_[43], _2059_[31], _2059_[22], _2059_[17], _2059_[5], _2059_[1:0] } = { _0992_, _0547_, _1282_, _1608_, _0822_, _1632_, _1474_, _1330_, _1382_, _1249_, _0697_, _0192_ };
  assign { _2060_[95:59], _2060_[50], _2060_[48:47], _2060_[45], _2060_[39:0] } = { _2033_[20:6], _0196_, _0325_, _2023_[13:12], _1469_, _1408_, _2023_[9:7], _0327_, _2023_[5:0], _0512_, _0023_, _0607_, _1625_, _0627_, _0099_, _0862_, _2057_[2:1], _1719_, _1393_, _1136_, _0306_, _0174_, _0657_, _1464_, _0359_, _0019_, _1368_, _1013_, _1266_, _0769_, _0997_, _0979_, _2001_[111], _1323_, _2001_[109], _1309_, _1081_, _2001_[106:103], _1351_, _2001_[101:99], _1353_, _2001_[97], _1359_, _0068_, _0671_, _1589_, _0191_, _1170_, _0003_, _1072_, _0438_, _1625_, _0290_ };
  assign _2061_[3] = _1554_;
  assign { _2062_[27], _2062_[20], _2062_[17], _2062_[5] } = { _0538_, _1849_, _1644_, _1642_ };
  assign { _2063_[42:41], _2063_[37:29], _2063_[27:0] } = { _1615_, _0147_, _1911_[14:8], _1284_, _0908_, _0059_, _0179_, _2042_[12:1], _1532_, _0419_, _0217_, _0220_, _0166_, _1343_, _1977_[25:24], _1243_, _1384_, _1669_, _0256_, _0617_, _0129_ };
  assign { _2064_[43:38], _2064_[36], _2064_[33:22], _2064_[13], _2064_[10:9], _2064_[6:0] } = { _1890_[11], _0350_, _0228_, _0177_, _0490_, _0552_, _1350_, _2024_[13:12], _1825_, _2024_[10:2], _1676_, _1049_, _1566_, _0408_, _0343_, _0627_, _1064_, _0572_, _0730_, _0505_ };
  assign { _2065_[39], _2065_[26] } = { _1400_, _1430_ };
  assign _2066_[5:2] = { _1937_, _1736_, _1480_ };
  assign { _2067_[5:3], _2067_[0] } = { _0926_, _0674_, _0610_, _0775_ };
  assign _2068_[30] = _1058_;
  assign { _2069_[22], _2069_[12:9], _2069_[7], _2069_[4:3], _2069_[1:0] } = { _1317_, _0202_, _0226_, _0531_, _1680_, _1458_, _0696_, _1649_, _0325_, _0922_ };
  assign { _2070_[17], _2070_[10], _2070_[4], _2070_[0] } = { _1201_, _1796_, _0165_, _0166_ };
  assign { _2071_[36], _2071_[21:14], _2071_[5] } = { _1824_, _1900_[86:79], _0427_ };
  assign _2072_[43:0] = { _1973_[25:24], _0504_, _1597_, _0684_, _1973_[20:19], _1970_[51:42], _1013_, _0662_, _0505_, _0277_, _2040_[20:11], _0618_, _1485_, _2040_[8], _1488_, _2040_[6:3], _1322_, _0661_, _1374_, _1035_, _0175_ };
  assign { _2073_[4], _2073_[2] } = { _0973_, _0280_ };
  assign _2074_[5:0] = { _2049_[83:82], _0246_, _0865_, _0354_, out_data[1920] };
  assign { _2075_[7], _2075_[5] } = { _0832_, _0927_ };
  assign _2076_[22] = _1610_;
  assign { _2077_[19], _2077_[14], _2077_[9], _2077_[6:4] } = { _1403_, _0742_, _0089_, _1227_, _1643_, _1542_ };
  assign { _2078_[15:14], _2078_[5] } = { _0579_, _1173_, _0826_ };
  assign _2079_[3:0] = { _0228_, _0613_, _0732_, _1015_ };
  assign { _2080_[22], _2080_[7], _2080_[3] } = { _0008_, _1707_, _0974_ };
  assign { _2081_[31:22], _2081_[20], _2081_[18], _2081_[15:0] } = { _1911_[14:8], _1284_, _0908_, _2063_[28], _1269_, _1376_, _0127_, _0337_, _0134_, _1633_, _0662_, _0988_, _0091_, _1627_, _0285_, _0999_, _1901_[66:63], _1575_, _1901_[61] };
  assign { _2082_[31], _2082_[26], _2082_[23], _2082_[18], _2082_[14:0] } = { _2035_[2], _0628_, _1223_, _1355_, _0025_, _0044_, _0149_, _0379_, _0607_, _1936_[47:44], _1612_, _1936_[42], _0418_, _1936_[40], _0619_, _0009_ };
  assign _2083_[6:0] = { _0361_, _0716_, _0163_, _0512_, _0681_, _1447_, _0198_ };
  assign { _2084_[6:2], _2084_[0] } = { _1906_[4:1], _0744_, _1420_ };
  assign _2085_[8:0] = { _2074_[6], _2049_[83:78], _0394_, _0650_ };
  assign _2086_[31:4] = { _1935_[79], _1157_, _1935_[77:72], _1953_[24:8], _1428_, _1953_[6], _1776_ };
  assign _2087_[30:0] = { _1966_[4], _0818_, _1966_[2], _0394_, _0092_, _0401_, _0140_, _1033_, _0228_, _2077_[20], _1403_, _2077_[18:15], _0742_, _2077_[13:10], _0089_, _2077_[8:7], _1227_, _1643_, _1542_, _2077_[3:0], _1689_ };
  assign _2088_[19] = _0577_;
  assign { _2089_[3], _2089_[1:0] } = { _1769_, _1526_, _0011_ };
  assign _2090_[10:7] = { _1945_[7:5], _1519_ };
  assign { _2091_[12], _2091_[10:0] } = { _0644_, _2014_[17:10], _1174_, _0550_, _0924_ };
  assign { _2092_[6], _2092_[4:0] } = { _1548_, _2064_[11], _1049_, _1566_, _2064_[8:7] };
  assign { _2093_[127], _2093_[76], _2093_[54:4] } = { _1071_, _1591_, _1899_[53:3] };
  assign { _2094_[102], _2094_[93], _2094_[68:56], _2094_[46], _2094_[44:29], _2094_[25], _2094_[23:21], _2094_[18], _2094_[13], _2094_[5], _2094_[2:0] } = { _1291_, _1263_, _0246_, _0332_, _0549_, _1195_, _0179_, _0183_, _0210_, _0303_, _0999_, _0598_, _0702_, _0612_, _0106_, _1732_, _1283_, _0103_, _2046_[6], _1756_, _2046_[4], _1094_, _2046_[2:0], _0043_, _0191_, _0151_, _1044_, _0704_, _0288_, _1021_, _1779_, _0691_, _1416_, _1781_, _0545_, _0346_, _1767_, _1645_, _0043_, _1799_ };
  assign { _2095_[126:118], _2095_[107:87], _2095_[39], _2095_[25], _2095_[23:22], _2095_[20:19], _2095_[11:0] } = { _2007_[8:1], _1441_, _1972_[25:23], _1686_, _0335_, _0076_, _1981_[11:9], _0299_, _0223_, _1981_[6:2], _1794_, _0189_, _0190_, _0694_, _0127_, _1516_, _1352_, _1661_, _1710_, _1162_, _1272_, _1585_, _0746_, _0466_, _0338_, _0784_, _0946_, _0703_, _1225_, _0619_, _0907_, _0419_, _0678_ };
  assign _2097_[4:0] = { _1037_, _1567_, _0299_, _0069_, _0032_ };
  assign { _2098_[39:19], _2098_[2:0] } = { _1984_[41:39], _1714_, _1984_[37:36], _0251_, _1984_[34:26], _1005_, _0057_, _1044_, _0808_, _1468_, _0289_, _0206_, _1392_ };
  assign { _2099_[8], _2099_[6] } = { _1840_, _1426_ };
  assign _2100_[27] = _0508_;
  assign { _2101_[162:116], _2101_[110:94], _2101_[89], _2101_[87:47], _2101_[39], _2101_[33], _2101_[26:0] } = { _2045_[8:5], _2012_[43:28], _1625_, _2012_[26:22], _1678_, _1222_, _2012_[19:2], _1613_, _1368_, _0566_, _1951_[123], _1122_, _1951_[121:119], _1609_, _0379_, _0096_, _1395_, _1380_, _0603_, _0152_, _0626_, _0683_, _1392_, _0910_, _1895_[35:26], _1111_, _1895_[24:20], _1757_, _1895_[18:3], _1634_, _0166_, _0752_, _1655_, _0198_, _0642_, _0438_, _0204_, _1163_, _1216_, _0658_, _1980_[23:6], _1367_, _1980_[4], _1681_, _1980_[2:0], _0518_, _0914_ };
  assign { _2102_[165:116], _2102_[52], _2102_[33], _2102_[12:0] } = { _0865_, _1651_, _0134_, _0289_, _0683_, _0681_, _0984_, _1247_, _0221_, _2096_, _0642_, _0399_, _1662_, _2073_[6:5], _0973_, _2073_[3], _0280_, _2073_[1:0], _0521_, _0692_, _0137_, _0681_, _0978_, _0631_ };
  assign _2104_[2:0] = { _0648_, _0354_, _1283_ };
  assign _2105_[37:0] = { _2035_[23:19], _1455_, _1507_, _2035_[16], _1674_, _2035_[14:2], _2082_[30:27], _0628_, _2082_[25:24], _1223_, _2082_[22:19], _1355_, _0265_, _1000_, _0238_ };
  assign { _2106_[24], _2106_[21] } = { _1728_, _0040_ };
  assign { _2107_[30:15], _2107_[12:3], _2107_[0] } = { _1995_[14], _0224_, _1995_[12], _1379_, _0041_, _2069_[8], _1458_, _2069_[6:5], _0696_, _1649_, _2069_[2], _0175_, _0176_, _1020_, _1601_, _2092_[14:7], _1548_, _2092_[5], _0368_ };
  assign { _2108_[84:81], _2108_[77], _2108_[75:46], _2108_[42:33], _2108_[30], _2108_[14:0] } = { _2011_[20:19], _0452_, _0182_, _1791_, _2053_[40:28], _1667_, _2053_[26:21], _1695_, _2053_[19:15], _1185_, _2053_[13:11], _0273_, _0217_, _0259_, _0657_, _1812_, _0984_, _0287_, _0020_, _0018_, _0510_, _1414_, _0031_, _0723_, _0453_, _0290_, _0144_, _0164_, _1043_, _1003_, _0076_, _0032_, _0712_, _0137_, _0581_, _0025_, _0274_ };
  assign _2109_[0] = _1546_;
  assign _2110_[45] = _1103_;
  assign { _2111_[51], _2111_[34], _2111_[28], _2111_[20], _2111_[3:0] } = { _1503_, _0661_, _2087_[31], _1200_, _0489_, _0469_, _1702_, _0866_ };
  assign { _2112_[94], _2112_[80:43], _2112_[27], _2112_[14], _2112_[11], _2112_[5] } = { _1803_, _2095_[130:127], _2007_[8:1], _1441_, _2095_[117:108], _1972_[25:22], _1687_, _1972_[20:11], _1666_, _0262_, _1604_, _0410_ };
  assign _2113_[10:0] = { out_data[544], _1933_[28:19] };
  assign _2114_[22:0] = { _0189_, _0759_, _1976_[19:16], _1335_, _1976_[14], _0172_, _0120_, _1568_, _1976_[10:9], _0604_, _1976_[7], _0945_, _1976_[5], _0602_, _1976_[3:0], _0857_ };
  assign { _2115_[7:5], _2115_[1] } = { _1479_, _1924_[7], _0847_, _0869_ };
  assign { _2116_[7], _2116_[4], _2116_[2] } = { _1499_, _1448_, _1523_ };
  assign { _2117_[5], _2117_[0] } = { _0432_, _0607_ };
  assign { _2119_[99:38], _2119_[29:28], _2119_[25], _2119_[19:18], _2119_[16], _2119_[13], _2119_[2:0] } = { _2038_[39:31], _0323_, _2080_[31:23], _0008_, _2080_[21:8], _1707_, _2080_[6:4], _0974_, _2080_[2:0], _0781_, _0559_, _0068_, _0059_, _1551_, _0228_, _0000_, _0857_, _1421_, _0265_, _0887_, _0113_, _0014_, _1704_, _0161_, _0671_, _0590_, _0217_, _0216_, _0605_, _1450_, _1638_, _1502_, _0828_, _2051_[9], _1106_, _1171_, _0030_, _0272_, _0631_ };
  assign { _2120_[99:33], _2120_[29], _2120_[15:0] } = { _1157_, _1935_[77:72], _1953_[24:8], _1428_, _1953_[6], _1776_, _0482_, _1761_, _1590_, _1929_[4:3], _1073_, _1627_, _1026_, _1409_, _2106_[30:25], _1728_, _2106_[23:22], _0040_, _2106_[20:0], _1762_, _0793_, _1425_, _1900_[72:70], _0389_, _1900_[68:66], _0833_, _1305_, _1900_[63], _0159_, _0466_, _0299_, _0924_ };
  assign { _2121_[97:44], _2121_[38:37], _2121_[34], _2121_[27], _2121_[21:2] } = { in_data[2137:2084], _0864_, _1346_, _1600_, _0653_, _2031_[66], _0328_, _2031_[64], _0007_, _1699_, _2031_[61:55], _1806_, _2031_[53], _0206_, _2031_[51], _1800_, _2031_[49:47] };
  assign _2122_[8:3] = { _1949_[9:5], _1273_ };
  assign _2123_[0] = _0129_;
  assign _2124_[8:0] = { _1452_, _1964_[75:74], _1647_, _1964_[72:68] };
  assign { _2125_[43], _2125_[12] } = { _0845_, _1277_ };
  assign { _2126_[48:45], _2126_[42:0] } = { _1699_, _2031_[61:59], _2101_[93:90], _0910_, _2101_[88], _1895_[35:26], _1111_, _1895_[24:20], _1757_, _1895_[18:3], _1027_, _0010_, _1554_, _1689_ };
  assign _2127_[1] = _1881_;
  assign _2128_[1] = _0782_;
  assign { _2130_[6], _2130_[3:1] } = { _1838_, _1492_, _1119_, _0952_ };
  assign _2132_[0] = _0282_;
  assign _2133_[0] = _1727_;
  assign { _2134_[5], _2134_[2:0] } = { _0003_, _0530_, _0018_, _0254_ };
  assign _2138_[35] = _1844_;
  assign { _2139_[72:67], _2139_[59], _2139_[54:53], _2139_[50], _2139_[48], _2139_[44], _2139_[42], _2139_[39:36], _2139_[31:30], _2139_[0] } = { _1901_[66:63], _1575_, _1901_[61], _1705_, _1743_, _0943_, _0345_, _1748_, _1837_, _1256_, _0337_, _1251_, _0590_, _0348_, _1354_, _1054_, _0277_ };
  assign _2140_[22:14] = { _1956_[30:24], _1618_, _1956_[22] };
  assign _2141_[18:0] = { _1901_[15:14], _0760_, _1901_[12:10], _0879_, _1901_[8:5], _1078_, _1901_[3], _0660_, _0311_, _1651_, _0057_, _0530_, _1017_ };
  assign { _2142_[84:81], _2142_[79:57], _2142_[55:54], _2142_[52:46], _2142_[42:41], _2142_[27], _2142_[17:5], _2142_[3:0] } = { _0447_, _0268_, _0991_, _0359_, _1134_, _1718_, _1422_, _0215_, out_data[416], _0529_, _0155_, _1974_[0], _2027_[10:9], _0889_, _2027_[7:5], _0260_, _2027_[3:1], _1107_, _0524_, _0299_, _0200_, _0296_, _0994_, _0702_, _0206_, _1164_, _1033_, _0314_, _0215_, _0978_, _0348_, _1830_, _0093_, _1775_, _2032_[66:54], _1304_, _0192_, _0164_, _0012_ };
  assign { _2143_[76], _2143_[2:0] } = { _1759_, _0228_, _0286_, _0692_ };
  assign { _2144_[63:56], _2144_[54:5] } = { _1891_[12:5], _1250_, _2072_[44], _1973_[25:24], _0504_, _1597_, _0684_, _1973_[20:19], _1970_[51:20], _1253_, _1970_[18:16], _1210_, _1682_, _1970_[13:11] };
  assign { _2145_[23:8], _2145_[6], _2145_[4], _2145_[0] } = { _1927_[19], _1565_, _1927_[17:6], _0853_, _0794_, _1062_, _1635_, _1093_ };
  assign { _2146_[20], _2146_[3:1] } = { _1763_, _0752_, _0519_, _0193_ };
  assign _2147_[4] = _1869_;
  assign { _2148_[49], _2148_[38], _2148_[29:28], _2148_[6] } = { _1851_, _0880_, _1934_[5:4], _1578_ };
  assign { _2149_[19:14], _2149_[7], _2149_[5:0] } = { _1063_, _0228_, _0680_, _0305_, _1064_, _0228_, _1152_, _0258_, _0297_, _1360_, _0132_, _0685_, _1363_ };
  assign _2150_[60:27] = _2143_[36:3];
  assign { _2151_[34:26], _2151_[24:5], _2151_[3:0] } = { _0918_, _0894_, _1838_, _2130_[5:4], _1492_, _1119_, _0952_, _2130_[0], _2146_[23:21], _1763_, _2146_[19:4], _1322_, _0075_, _0678_, _1245_ };
  assign _2153_[23] = _1508_;
  assign { _2154_[34], _2154_[31:0] } = { _1080_, _1338_, _0851_, _0242_, _0540_, _0318_, _0417_, _2044_[8:6], _0668_, _2044_[4:1], _1461_, _0905_, _0323_, _0076_, _1941_[13:1], _0895_ };
  assign _2155_[1] = _1871_;
  assign { _2158_[47], _2158_[39], _2158_[33] } = { _1300_, _1563_, _1489_ };
  assign { _2159_[47:8], _2159_[1] } = { _1907_[55:25], _1535_, _1907_[23:16], _1842_ };
  assign _2160_[23:0] = { _0749_, _0590_, _1901_[66:63], _1575_, _1901_[61], _0855_, _1459_, _0058_, _0298_, _1936_[47:44], _1612_, _1936_[42], _0418_, _1936_[40], _1121_, _0366_, _0548_, _0649_ };
  assign _2161_[28:12] = { _1901_[15:14], _0760_, _1901_[12:10], _0879_, _1901_[8:5], _1078_, _1901_[3], _0711_, _0600_, _0503_, _0524_ };
  assign { _2162_[17], _2162_[15], _2162_[8] } = { _0874_, _1766_, _1155_ };
  assign _2163_[24:0] = { _0228_, _1228_, _0748_, _1655_, _1051_, _0703_, _1088_, _1348_, _0566_, _0358_, _0936_, _0221_, _1090_, _0323_, _1951_[123], _1122_, _1951_[121:119], _1609_, _0267_, _0899_, _0279_, _0034_, _0988_ };
  assign { _2164_[23], _2164_[19:17], _2164_[11:3] } = { _0601_, _1997_, _2154_[39:35], _1080_, _2154_[33:32], _1338_ };
  assign { _2165_[46:12], _2165_[10:0] } = { _2100_[161:152], _1663_, _0288_, _0844_, _1713_, _0835_, _1808_, _0216_, _1038_, _1254_, _0468_, _2006_[6], _0404_, _2006_[4:3], _1931_[3], _1308_, _0513_, _1095_, _1023_, _2147_[5], _1869_, _2147_[3:0], _1187_, _0626_, _0678_, _0682_, _0436_, _0659_, _0502_, _0178_, _1377_, _0642_, _0303_ };
  assign { _2166_[45], _2166_[35:14], _2166_[12:0] } = { _1100_, _0548_, _2015_[20:2], _1369_, _2015_[0], _1609_, _2027_[10:9], _0889_, _2027_[7:5], _0260_, _2027_[3:1], _1107_, _0464_ };
  assign _2167_[5] = _1524_;
  assign { _2168_[165], _2168_[110:57] } = { _1521_, _1989_[54:33], _1344_, _1989_[31:5], _1792_, _1989_[3:2], _1992_[8] };
  assign { _2169_[169:102], _2169_[100:57], _2169_[54], _2169_[44], _2169_[39], _2169_[34:0] } = { _1972_[13:11], _2112_[42:28], _1666_, _2112_[26:15], _0262_, _2112_[13:12], _1604_, _2112_[10:6], _0410_, _2112_[4:1], _1203_, _0189_, _0228_, _0189_, _1153_, _1893_[10:7], _1034_, _1893_[5:4], _1374_, _1787_, _0126_, _1328_, _0287_, _0238_, _0134_, _0304_, _0205_, _0096_, _0200_, _2105_[43:38], _2035_[23:19], _1455_, _1507_, _2035_[16], _1674_, _2035_[14:2], _2082_[30:27], _0628_, _2082_[25:24], _1223_, _2082_[22:19], _1355_, _2082_[17:15], _0451_, _1793_, _1324_, _2000_[59:50], _1570_, _2000_[48:46], _1314_, _1419_, _0391_, _2000_[42:35], _1747_, _2000_[33:31], _1307_, _2000_[29:27], _1318_, _0106_ };
  assign { _2170_[169:85], _2170_[69:38], _2170_[30], _2170_[25], _2170_[8], _2170_[3:0] } = { _2000_[122:108], _1361_, _2000_[106:100], _1506_, _2000_[98], _0113_, _2000_[96:92], _0313_, _2000_[90:86], _0737_, _2000_[84:83], _0237_, _1206_, _0573_, _1046_, _0084_, _0270_, _0464_, _0638_, _0272_, _0356_, _0232_, _1283_, _0071_, _2164_[29:24], _0601_, _2164_[22:20], _1997_, _2164_[16:12], _2154_[39:35], _1080_, _2154_[33:32], _1338_, _2164_[2:0], _0194_, _0317_, _2070_[32:18], _1201_, _2070_[16:11], _1796_, _2070_[9:5], _0165_, _2070_[3:1], _1008_, _1332_, _0169_, _1203_, _0354_, _0232_, _0241_ };
  assign { _2173_[20], _2173_[2:0] } = { _1460_, _0163_, _1443_, _1471_ };
  assign { _2174_[8:6], _2174_[1] } = { _0444_, _1572_, _1653_, _0969_ };
  assign { _2175_[6], _2175_[3:2] } = { _1252_, _0839_, _0836_ };
  assign { _2177_[33:18], _2177_[14], _2177_[4] } = { _2172_[16:2], _0009_, _1495_, _1191_ };
  assign { _2178_[78:43], _2178_[25], _2178_[17:10], _2178_[5:3], _2178_[1:0] } = { _1903_[38:36], _1213_, _1903_[34:5], _0645_, _0009_, _0396_, _1203_, _1301_, _0071_, _0587_, _1539_, _1935_[26:25], _0481_, _0217_, _0603_, _1046_, _0724_, _0672_ };
  assign _2181_[1] = _0228_;
  assign { _2182_[76:53], _2182_[42], _2182_[25] } = { _1925_[30:7], _0584_, _0976_ };
  assign { _2183_[49], _2183_[28:13], _2183_[8], _2183_[2:0] } = { _1349_, _2079_[21:16], _0571_, _1977_[25:24], _1243_, _1384_, _1669_, _0256_, _0041_, _1720_, _0656_, _0906_, _0044_, _0888_, _0367_ };
  assign { _2184_[12], _2184_[5] } = { _1630_, _1740_ };
  assign { _2185_[64:59], _2185_[57], _2185_[31:23], _2185_[5] } = { _2139_[61:60], _1705_, _2139_[58:56], _0116_, _2176_, _1475_, _1703_ };
  assign { _2186_[28:5], _2186_[1:0] } = { _1952_[56:45], _1232_, _1494_, _1952_[42], _0803_, _1952_[40:33], _0932_, _1298_ };
  assign { _2187_[22:9], _2187_[3] } = { _1941_[37:24], _1745_ };
  assign { _2188_[18], _2188_[4:0] } = { _0459_, _0352_, _1691_, _0176_, _1422_, _0796_ };
  assign { _2189_[71:69], _2189_[43], _2189_[36], _2189_[33] } = { _1923_[7:5], _1641_, _1159_, _1588_ };
  assign { _2190_[78:75], _2190_[73:0] } = { _1144_, _0289_, _1579_, _1573_, _0071_, _1478_, out_data[1184], _0560_, _1129_, _0565_, _0599_, _0206_, _0754_, _0529_, _1009_, _0043_, _1102_, _0633_, _0162_, _1959_[7], _1202_, _2116_[8], _1499_, _2116_[6:5], _1448_, _2116_[3], _1523_, _2116_[1:0], _0325_, _1425_, _1286_, _0511_, _0872_, _2174_[9], _0444_, _1572_, _1653_, _2174_[5:2], _0969_, _2174_[0], _0343_, _0285_, _1614_, _0695_, _0019_, _1348_, _2077_[20], _1403_, _2077_[18:15], _0742_, _2077_[13:10], _0089_, _2077_[8:7], _1227_, _1643_, _1542_, _2077_[3:0], _0893_, _0420_, _1235_, _0157_, _0358_, _0654_ };
  assign _2191_[6:0] = _1914_[46:40];
  assign _2192_[13] = _1944_[35];
  assign { _2194_[10], _2194_[8:5], _2194_[3:0] } = { _0726_, _2134_[6], _0003_, _2134_[4:3], _0503_, _2165_[11], _1187_, _0004_ };
  assign _2195_[5:0] = { _0412_, _1827_, _1625_, _1610_, _0649_, _0047_ };
  assign _2196_[60] = _1861_;
  assign { _2197_[154:92], _2197_[89], _2197_[81:78], _2197_[25:0] } = { _1971_[24:19], _0922_, _1971_[17:13], _1525_, _1971_[11:3], _0228_, _0285_, _0179_, _0317_, _0631_, _0157_, _1554_, _1468_, _2098_[18:3], _1208_, _1174_, _0704_, _1828_, _0701_, _0298_, _0817_, _0609_, _1017_, _0848_, _0012_, _0009_, _0756_, _0193_, _0217_, _0014_, _0627_, _0877_, _0271_, _0032_, _1481_, _1835_, _0467_, _0337_, _1170_, _1561_, _1456_, _1447_, _1554_, _0669_, _1374_, _0237_, _2152_, _0812_, _1203_, _0368_, _0103_, _0478_, _0027_, _0115_, _0343_, _1585_, _0987_, _1552_, _0709_ };
  assign _2198_[5] = _1545_;
  assign { _2199_[47:28], _2199_[20], _2199_[15:0] } = { _2183_[78:59], _0996_, _2010_[3:1], _0240_, _0844_, _1713_, _1433_, _0251_, _2193_ };
  assign { _2200_[41:40], _2200_[19:0] } = { _1855_, _0923_, _0202_, _1394_, _1046_, _1270_, _0807_, _1154_, _0609_, _2127_[6:2], _1881_, _2127_[0], _0217_, _0670_, _1615_, _0381_, _0347_, _0799_ };
  assign { _2201_[11:6], _2201_[4:0] } = { _0289_, _0005_, _0633_, _0162_, _1959_[7], _1202_, _1095_, _1689_, _0891_, _0848_, _0638_ };
  assign { _2202_[3:2], _2202_[0] } = { _1184_, _1773_, _1774_ };
  assign { _2203_[17], _2203_[9], _2203_[7:3] } = { _1671_, _1571_, _1938_[8:5], _0131_ };
  assign _2204_[1:0] = { _1672_, _0821_ };
  assign { _2205_[17:10], _2205_[2] } = { _0726_, _2194_[9], _2134_[6], _0003_, _2134_[4:3], _2194_[4], _1091_, _1693_ };
  assign _2206_[6] = _0981_;
  assign _2208_[0] = _1281_;
  assign { _2209_[31:30], _2209_[15], _2209_[13:0] } = { _0972_, _2201_[12], _1620_, _1966_[77:67], _0179_, _0284_, _0116_ };
  assign _2210_[3] = _1875_;
  assign { _2211_[6], _2211_[2:0] } = { _1541_, _0146_, _1121_, _0687_ };
  assign { _2213_[17:4], _2213_[2:0] } = { _0208_, _1114_, _1270_, _0192_, _0159_, _1636_, _2117_[8:6], _0432_, _2117_[4:1], _0347_, _0421_, _1135_ };
  assign { _2214_[23], _2214_[21:0] } = { _1490_, _0034_, _0238_, _2139_[66:60], _1705_, _2139_[58:55], _1743_, _0943_, _2139_[52:51], _0507_, _1139_, _1072_, _1551_ };
  assign _2215_[1:0] = { _1559_, _2213_[23] };
  assign { _2216_[98], _2216_[85], _2216_[79], _2216_[61:3], _2216_[0] } = { _1511_, _0734_, _1278_, _1952_[215:214], _1083_, _1952_[212:206], _1246_, _1952_[204:184], _1389_, _1952_[182:177], _0344_, _1952_[175:165], _1194_, _1952_[163:157], _0635_ };
  assign { _2217_[41:25], _2217_[20] } = { _1904_[38:22], _1226_ };
  assign { _2218_[43:13], _2218_[0] } = { _1942_[86:58], _0905_, _1170_, _0563_ };
  assign { _2219_[30:10], _2219_[7:0] } = { _2069_[32:23], _1317_, _2069_[21:18], _0545_, _0796_, _0258_, _0232_, _0415_, _1558_, _0284_, _0449_, _1233_, _0021_, _0134_, _0324_, _0165_, _1371_ };
  assign { _2220_[82:76], _2220_[14], _2220_[11:0] } = { _2093_[75:71], _0271_, _0619_, _1032_, out_data[1344], _1254_, _0468_, _2006_[6], _0404_, _2006_[4:3], _1931_[3], _1308_, _0513_, _0710_, _0827_ };
  assign { _2221_[82:77], _2221_[74], _2221_[70:68], _2221_[58], _2221_[55:53], _2221_[51:49], _2221_[47:36], _2221_[9:0] } = { _2090_[12:11], _1945_[7:6], _0475_, _0166_, _0536_, _1688_, _1815_, _1432_, _1543_, _0164_, _1019_, _0342_, _0766_, _0415_, _0663_, _0221_, _0176_, _1233_, _1031_, _1134_, _1436_, _0562_, _0369_, _1805_, _2009_[2], _0819_, _1807_, _1956_[18:15], _0506_, _1956_[13:12], _0651_, _0250_, _1641_ };
  assign { _2223_[42:16], _2223_[1:0] } = { _1896_[35:24], _1594_, _1896_[22:12], _1712_, _1896_[10:9], _0733_, _1110_ };
  assign _2224_[15] = _0916_;
  assign { _2225_[64:63], _2225_[60:58], _2225_[56:11], _2225_[9], _2225_[3:2], _2225_[0] } = { _2006_[3], _1931_[3], _0464_, _0893_, _1809_, _1633_, _0808_, _2142_[45:43], _1830_, _0093_, _2142_[40:28], _1775_, _2142_[26:18], _2032_[66:54], _2142_[4], _1239_, _1866_, _0962_, _0971_, _0216_, _0092_ };
  assign { _2226_[67:34], _2226_[23:0] } = { _2112_[85:81], _2095_[130:127], _2007_[8:1], _1441_, _2095_[117:111], _1396_, _1131_, _0217_, _0228_, _0022_, _0469_, _1089_, _0164_, _0471_, _1921_, _0530_, _0456_, _0612_, _1225_, _2177_[17:15], _1495_, _2177_[13:5], _1191_, _2177_[3:0], _0302_ };
  assign { _2227_[38:36], _2227_[34:23], _2227_[11:1] } = { _2155_[4:2], _0572_, _0472_, _0825_, _0694_, _0712_, _0598_, _0367_, _0807_, _0710_, _0016_, _0715_, _0490_, _2211_[13:7], _1541_, _2211_[5:3] };
  assign { _2228_[47], _2228_[40:33], _2228_[26] } = { _0541_, _1894_[55:48], _1262_ };
  assign { _2229_[67:38], _2229_[30:26], _2229_[24:0] } = { _2014_[16:10], _1988_[54:51], _0291_, _1988_[49], _1383_, _1988_[47:46], _1697_, _1988_[44], _1153_, _1893_[10:7], _1034_, _1893_[5:4], _1374_, _1787_, _0126_, _1328_, _0867_, _0641_, _1752_, _1721_, _1836_, _0548_, _2015_[20:2], _1369_, _2015_[0], _0799_, _0004_, _1760_ };
  assign _2230_[8] = _0078_;
  assign { _2231_[197:160], _2231_[158], _2231_[155:154], _2231_[152], _2231_[150:95], _2231_[80:53], _2231_[44:3], _2231_[0] } = { _2117_[7:6], _0432_, _2117_[4:1], _2213_[3], _0453_, _1470_, _0132_, _2008_[14:3], _1531_, _1068_, _2008_[0], _0094_, _0101_, _2127_[6:2], _1881_, _2127_[0], _1501_, _1846_, _1248_, _0045_, _1751_, _1536_, _0216_, _0221_, _1112_, _1530_, _0588_, _1890_[11], _0350_, _0716_, _1890_[8:6], _0294_, _2157_, _0321_, _0106_, _0289_, _0704_, _2165_[11], _1187_, _2200_[47:42], _1855_, _0923_, _2200_[39:20], _1988_[41:38], _0130_, _1988_[36], _0725_, _1988_[34:27], _1406_, _1175_, _1988_[24], _0921_, _1988_[22], _1819_, _1988_[20:19], _0778_, _0059_, _0703_, _2050_[9:5], _1164_, _2050_[3:2], _1296_, _2050_[0], _0682_, _0069_, _0590_, _0315_, _0671_, _0484_, _0419_ };
  assign { _2232_[7], _2232_[4], _2232_[2:0] } = { _0063_, _0375_, _1544_, _1691_, _0899_ };
  assign _2233_[0] = _0965_;
  assign { _2234_[32:22], _2234_[5:4], _2234_[2:1] } = { _2001_[123:113], _2132_[1], _0791_, _0423_, _0193_ };
  assign { _2235_[45:35], _2235_[21] } = { _0516_, _1958_[13:4], _0006_ };
  assign { _2236_[66:40], _2236_[31], _2236_[24:23], _2236_[18:6], _2236_[3:0] } = { _2153_[25:24], _1508_, _2153_[22:0], _1005_, _1700_, _1224_, _0664_, _2215_[7:2], _1559_, _2213_[23:18], _2208_[3:1], _1281_ };
  assign { _2237_[40:32], _2237_[28] } = { _0986_, _1908_[14:13], _1564_, _1908_[11:10], _0535_, _1908_[8], _0814_, _1219_ };
  assign { _2238_[86], _2238_[80:74], _2238_[71], _2238_[56:40], _2238_[30:7], _2238_[4] } = { _1522_, _2212_, _0378_, _1673_, _2016_[21:6], _1943_[111], _1768_, _1943_[109:89], _1007_, _1771_ };
  assign { _2240_[72:34], _2240_[32:10] } = { _2062_[41:28], _0538_, _2062_[26:21], _1849_, _2062_[19:18], _1644_, _2062_[16:6], _1642_, _2062_[4], _1463_, _2063_[43], _1615_, _0147_, _2063_[40:38], _1911_[14:8], _1284_, _0908_, _2063_[28], _2081_[21], _1269_, _2081_[19], _1376_, _2081_[17:16], _0642_ };
  assign { _2241_[38:14], _2241_[3:2] } = { _1936_[79:55], _1742_, _1686_ };
  assign { _2242_[20], _2242_[17], _2242_[15], _2242_[0] } = { _1316_, _0616_, _1378_, _1778_ };
  assign _2243_[8:0] = { _0768_, _0276_, _0116_, _0127_, _1046_, _0626_, _0227_, _1229_, _1518_ };
  assign { _2244_[80], _2244_[66], _2244_[55:4] } = { _0970_, _1319_, _2059_[95:89], _0992_, _2059_[87:76], _0547_, _2059_[74:71], _1282_, _2059_[69:67], _1608_, _2059_[65:55], _0822_, _2059_[53:44] };
  assign { _2245_[82:80], _2245_[78:73], _2245_[69:38], _2245_[33:31], _2245_[27:0] } = { _0049_, _0752_, _1070_, _1313_, _0624_, _2141_[22:19], _1984_[46:39], _1714_, _1984_[37:36], _0251_, _1984_[34:15], _1922_, _2091_[14:13], _0644_, _2091_[11], _2014_[17:10], _1988_[54:51], _0291_, _1988_[49], _1383_, _1988_[47:46], _1697_, _1988_[44:43], _0228_, _0191_, _0325_, _0453_ };
  assign _2246_[1] = _0086_;
  assign { _2248_[6], _2248_[3:0] } = { _1827_, _0217_, _1024_, _2222_ };
  assign { _2249_[26:25], _2249_[6:0] } = { _1652_, _1241_, _0324_, _1148_, _0590_, _0228_, _0138_, _0587_, _0182_ };
  assign { _2250_[41], _2250_[20:1] } = { _1749_, _2128_[16:2], _0782_, _2128_[0], _1017_, _0044_, _0733_ };
  assign { _2251_[14:13], _2251_[0] } = { _1490_, _2214_[22], _0924_ };
  assign _2253_[4:3] = { _0678_, _0335_ };
  assign { _2254_[52], _2254_[50:19], _2254_[17], _2254_[13], _2254_[11], _2254_[1] } = { _0878_, _2054_[40:39], _2039_[13:11], _1417_, _2054_[34:31], _1683_, _2054_[29:19], _1538_, _2054_[17:16], _1029_, _2054_[14:9], _1717_, _1404_, _1798_, _0167_ };
  assign _2255_[31:0] = out_data[1503:1472];
  assign _2256_[48:5] = { _1969_[51:36], _0677_, _1969_[34:29], _0985_, _1969_[27:8] };
  assign _2257_[35:4] = out_data[63:32];
  assign _2258_[59:15] = { _2001_[139:138], _0211_, _2001_[136:113], _2234_[21:6], _2132_[1], _0791_ };
  assign { _2259_[53:21], _2259_[18:1] } = { _2219_[43:31], _2069_[32:23], _1317_, _2069_[21:13], _2085_[9], _2074_[6], _2049_[83:72], _1121_, _2049_[70:69], _1670_ };
  assign { _2260_[22:20], _2260_[12] } = { _2056_[3:1], _0806_ };
  assign { _2261_[103], _2261_[67:31], _2261_[25] } = { _1104_, _2026_[43:34], _0842_, _2026_[32:11], _1097_, _2026_[9:7], _1045_ };
  assign { _2262_[109:57], _2262_[53], _2262_[51:0] } = { _0597_, _2048_[51:50], _1423_, _2048_[48:47], _2005_[10:8], _1327_, _2005_[6:4], _2048_[39:38], _1150_, _2048_[36], _1010_, _2048_[34:28], _0477_, _0651_, _0163_, _1203_, _0522_, _1206_, _1113_, _0408_, _0811_, _1956_[18:15], _0506_, _1956_[13:12], _0591_, _0795_, _0275_, _0887_, _0110_, _0334_, _0926_, _0674_, _0610_, _2067_[2:1], _0775_, _1690_, _2025_[43:40], _1785_, _2025_[38:34], _1510_, _2025_[32:27], _0896_, _2025_[25], _1556_, _0114_, _0319_, _2041_[32:31], _1755_, _2041_[29:24], _0233_, _0499_, _2114_[25:23], _0071_, _1964_[67], _0364_, _1888_[13], _0036_, _0706_, _1888_[10:5], _0673_, _1964_[55], _1679_, _1311_ };
  assign _2263_[59:5] = { _2101_[165:163], _2045_[8:5], _2012_[43:28], _1625_, _2012_[26:22], _1678_, _1222_, _2012_[19:2], _1613_, _2101_[115:111] };
  assign { _2264_[90:74], _2264_[58], _2264_[51], _2264_[16:6] } = { _1503_, _2111_[50:35], _0968_, _1802_, _2043_[12:2] };
  assign { _2265_[47], _2265_[37:2] } = { _1333_, _2241_[39], _1936_[79:55], _2241_[13:4] };
  assign _2266_[95:4] = { _2183_[102:50], _1349_, _2183_[48:29], _2079_[21:4] };
  assign _2267_[6] = _1214_;
  assign { _2268_[77:44], _2268_[37:3] } = { _1961_[34:1], _2038_[80:48], _1039_, _2038_[46] };
  assign { _2269_[11], _2269_[7:5] } = { _0892_, _1050_, _0329_, _1813_ };
  assign _2270_[66:4] = { _0667_, _2094_[130:103], _1291_, _2094_[101:94], _1263_, _2094_[92:69] };
  assign _2271_[37] = _1694_;
  assign { _2272_[14], _2272_[12:9] } = { _2252_, _2104_[6:3] };
  assign _2273_[27:1] = { _1919_[31:17], _0557_, _1919_[15:7], _1882_, _1919_[5] };
  assign _2274_[31:0] = { _2209_[32], _0972_, _2201_[12], _2209_[29:16], _1620_, _2209_[14], _1966_[77:65] };
  assign { _2276_[51], _2276_[39:18], _2276_[14] } = { _1637_, _2123_[22:1], _1860_ };
  assign { _2278_[56], _2278_[35], _2278_[31] } = { _1886_[16], _1738_, out_data[1600] };
  assign { _2279_[41:20], _2279_[4] } = { _2083_[28:7], _0556_ };
  assign { _2280_[58], _2280_[30] } = { _1482_, _0903_ };
  assign { _2281_[64], _2281_[55], _2281_[50:33] } = { _1280_, _1583_, _2163_[42:25] };
  assign { _2282_[101], _2282_[98:72], _2282_[59:19], _2282_[10] } = { _0938_, _2160_[50:24], _2149_[60:20], _1444_ };
  assign { _2283_[85], _2283_[69:53], _2283_[17] } = { _1240_, _2129_, _0365_ };
  assign { _2284_[39], _2284_[31], _2284_[6] } = { _1477_, _1143_, _1437_ };
  assign { _2285_[75], _2285_[70], _2285_[54:26] } = { _1398_, _1611_, _2248_[35:7] };
  assign { _2286_[8], _2286_[5] } = { _0966_, _1146_ };
  assign { _2287_[25], _2287_[22], _2287_[15:9] } = { _0500_, _0720_, _2180_ };
  assign { _2288_[3], _2288_[1] } = { _0491_, _1622_ };
  assign _2289_[120:12] = { _2143_[84:77], _1759_, _2143_[75:3], _2150_[26:0] };
  assign _2290_[45:11] = _2097_[39:5];
  assign _2291_[10] = _1628_;
  assign _2292_[1] = _1709_;
  assign _2293_[12:2] = { _2166_[46], _1100_, _2166_[44:36] };
  assign { _2294_[5], _2294_[3] } = { _0520_, _1140_ };
  assign { _2295_[27], _2295_[11] } = { _0002_, _0750_ };
  assign { _2296_[6], _2296_[3] } = { _1581_, _0388_ };
  assign _2297_[2] = _1735_;
  assign _2298_[29:1] = { _1954_[28:12], _1872_, _1954_[10:9], out_data[1952], _1954_[7:0] };
  assign _2299_[8] = _1271_;
  assign _2300_[14] = _1730_;
  assign _2301_[22:2] = { _2173_[23:21], _1460_, _2173_[19:3] };
  assign _2302_[52:2] = { _2159_[50:48], _1907_[55:25], _1535_, _1907_[23:16], _2159_[7:2], _1842_, _2159_[0] };
  assign _2303_[6] = _1859_;
  assign _2305_[26:11] = { _2251_[16:15], _1490_, _2214_[22], _2251_[12:1] };
  assign _2306_[25] = _1854_;
  assign { _2307_[23], _2307_[21], _2307_[9] } = { _1576_, _0428_, _1856_ };
  assign _2308_[99:61] = { _2178_[81:79], _1903_[38:36], _1213_, _1903_[34:3] };
  assign { _2309_[6], _2309_[4] } = { _1874_, _1180_ };
  assign { _2310_[49:45], _2310_[13:4] } = { _2195_[10:6], _2181_[11:2] };
  assign { _2311_[47], _2311_[15] } = { _0863_, _1623_ };
  assign _2312_[0] = _0474_;
  assign _2313_[21] = _1782_;
  assign { _2314_[21:17], _2314_[5] } = { _1946_[13:9], _2239_ };
  assign { _2315_[72], _2315_[27] } = { _1584_, _2247_ };
  assign { _2316_[5], _2316_[1] } = { _1582_, _1605_ };
  assign _2317_[42:5] = { _2250_[70:42], _1749_, _2250_[40:33] };
  assign { _2318_[6:5], _2318_[3] } = { _2253_[6:5], _1877_ };
  assign _2319_[34:31] = _2243_[12:9];
  assign _2320_[11] = _0583_;
  assign { _2321_[51:35], _2321_[16], _2321_[14], _2321_[0] } = { _1909_[39:35], _0254_, _1909_[33:25], _2204_[2], _1672_, _1848_, _1789_, _2277_ };
  assign { _2322_[56], _2322_[37:4] } = { _0073_, _2249_[40:27], _1652_, _1241_, _2249_[24:7] };
  assign { _2323_[33:24], _2323_[15] } = { _1948_, _1297_ };
  assign out_data[224] = out_data[256];
endmodule
